netcdf line_z_cra {
dimensions:
	instance = 2 ;
	node = 5 ;
variables:
	int geometry_container ;
		geometry_container:geometry_type = "line" ;
		geometry_container:node_coordinates = "x y z" ;
		geometry_container:node_count = "node_count" ;
	double x(node) ;
		x:axis = "X" ;
	double y(node) ;
		y:axis = "Y" ;
	double z(node) ;
		z:axis = "Z" ;
	int node_count(instance) ;
		node_count:long_name = "count of coordinates in each instance geometry" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 geometry_container = _ ;

 x = 3, 1, 4, 7, 8 ;

 y = 1, 3, 4, 9, 10 ;

 z = NaN, NaN, NaN, 90, 100 ;

 node_count = 3, 2 ;
}
