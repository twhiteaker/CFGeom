netcdf polygon_hole_cra {
dimensions:
	instance = 2 ;
	node = 10 ;
	part = 3 ;
variables:
	int geometry_container ;
		geometry_container:geometry_type = "polygon" ;
		geometry_container:node_coordinates = "x y" ;
		geometry_container:node_count = "node_count" ;
		geometry_container:part_node_count = "part_node_count" ;
		geometry_container:interior_ring = "interior_ring" ;
	double x(node) ;
		x:axis = "X" ;
	double y(node) ;
		y:axis = "Y" ;
	int node_count(instance) ;
		node_count:long_name = "count of coordinates in each instance geometry" ;
	int part_node_count(part) ;
		part_node_count:long_name = "count of nodes in each geometry part" ;
	int interior_ring(part) ;
		interior_ring:long_name = "type of each polygon geometry part" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 geometry_container = _ ;

 x = 10, 5, 0, 1, 5, 9, 20, 15, 11, 15 ;

 y = 0, 5, 0, 1, 4, 1, 20, 25, 20, 15 ;

 node_count = 6, 4 ;

 part_node_count = 3, 3, 4 ;

 interior_ring = 0, 1, 0 ;
}
