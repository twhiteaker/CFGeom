netcdf multipoint_vlen {
types:
  double(*) node_VLType ;
dimensions:
	instance = 2 ;
variables:
	int geometry_container ;
		geometry_container:geometry_type = "point" ;
		geometry_container:node_coordinates = "x y" ;
	node_VLType x(instance) ;
		x:axis = "X" ;
	node_VLType y(instance) ;
		y:axis = "Y" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 geometry_container = _ ;

 x = {1}, {1, 4} ;

 y = {1}, {4, 3} ;
}
