netcdf nwm_bullcreek {
  dimensions:
    time = 15;
    station = 20;
  variables:
    int time(time);
      time:long_name = "time";
      time:standard_name = "time";
      time:units = "seconds since 2016-11-07 20:00 UTC";

    int station_id(station);
      station_id:long_name = "Station id";

    float streamflow(time, station);
      streamflow:long_name = "River Flow";
      streamflow:units = "meter^3 / sec";

  // global attributes:
  :Conventions = "Unidata Observation Dataset v1.0";
  :cdm_datatype = "Station";
  :model_initialization_time = "2016-11-07_19:00:00";
  :station_dimension = "station";
  :missing_value = -8.9999998E15f; // float
  :stream_order_output = 1; // int
  :model_output_valid_time = "2016-11-08_04:00:00";

 data:
time =
  0, 3600, 7200, 10800, 14400, 18000, 21600, 25200, 28800, 32400, 36000, 39600, 43200, 46800, 50400 ;
station_id =
  5781157, 5781193, 5781183, 5781189, 5781173, 5781133, 5781163, 5781131, 5781141, 5781171, 5781159, 5781129, 5781139, 5781149, 5781185, 5781187, 5781145, 5781781, 5781191, 5781811 ;
streamflow =
    0.01282661, 0.42142317, 0.6132626, 0.36973292, 0.27779508, 0.07792676, 0.21289445, 0.022072816, 0.02037233, 0.29445773, 0.054952983, 0.055809632, 0.0016493346, 0.0068484014, 0.010602541, 0.022358151, 0.007151061, 0.0069096438, 0.04669686, -8.9999998E15,
    0.0128412, 0.30901003, 0.2857758, 0.27685326, 0.17878114, 0.07953472, 0.14906085, 0.022236675, 0.020542009, 0.10206464, 0.028738864, 0.05726831, 0.0016436642, 0.007000346, 0.010707803, 0.0057302667, 0.0073062116, 0.0070617246, 0.03053636, -8.9999998E15,
    0.012942635, 0.2950936, 0.2652008, 0.2710669, 0.17189544, 0.07931047, 0.13895877, 0.022362068, 0.02085562, 0.09134504, 0.032691292, 0.0569133, 0.0014596866, 0.0072410507, 0.010852132, 0.008282697, 0.0075517693, 0.0073028416, 0.023084112, -8.9999998E15,
    0.013025638, 0.2963086, 0.2631511, 0.27260152, 0.16236217, 0.0797341, 0.14336994, 0.022470536, 0.020963334, 0.09949419, 0.018426947, 0.05722875, 0.0014604526, 0.0072657303, 0.010920734, 0.008298121, 0.007576539, 0.0073275077, 0.023205092, -8.9999998E15,
    0.013108982, 0.30076107, 0.26495057, 0.27668196, 0.16340037, 0.08016156, 0.1442623, 0.02257986, 0.02107178, 0.10008767, 0.018518273, 0.0575469, 0.0014613364, 0.0072907805, 0.010989491, 0.008349704, 0.0076017086, 0.0073525496, 0.023355357, -8.9999998E15,
    0.013192658, 0.30424386, 0.26669532, 0.27994442, 0.16430004, 0.08059214, 0.145032, 0.022689886, 0.021180851, 0.10092157, 0.01864383, 0.057867453, 0.0014622996, 0.007316067, 0.011058502, 0.0084016435, 0.0076271477, 0.007377835, 0.023506908, -8.9999998E15,
    0.0132764615, 0.31614244, 0.27220803, 0.28619307, 0.16763578, 0.081025265, 0.1481796, 0.0228003, 0.021290282, 0.1030719, 0.01877265, 0.058190178, 0.0014632859, 0.007341582, 0.011501618, 0.013693551, 0.007652818, 0.0074033495, 0.029268358, -8.9999998E15,
    0.013360315, 0.31056792, 0.27054676, 0.28572553, 0.16622692, 0.08146068, 0.14667702, 0.022910941, 0.021399913, 0.10272537, 0.018904794, 0.058514945, 0.0014642992, 0.0073672463, 0.011192806, 0.00850965, 0.0076786387, 0.0074290126, 0.023817388, -8.9999998E15,
    0.013444155, 0.31257704, 0.27211815, 0.28770262, 0.16698666, 0.08189801, 0.14738096, 0.023021765, 0.021509703, 0.10362644, 0.019040179, 0.058841452, 0.0014653369, 0.007393077, 0.011266076, 0.0085587995, 0.0077046314, 0.0074548433, 0.023966836, -8.9999998E15,
    0.013527915, 0.31500065, 0.27398166, 0.2899553, 0.16798826, 0.08233685, 0.14817467, 0.023132667, 0.021619545, 0.10449046, 0.019178566, 0.059169404, 0.0014664014, 0.007419034, 0.011335222, 0.008611545, 0.00773075, 0.0074808, 0.024121437, -8.9999998E15,
    0.013611533, 0.40163192, 0.3468528, 0.36964124, 0.17151178, 0.08277698, 0.14897789, 0.023243539, 0.021729335, 0.16329302, 0.019319706, 0.05949866, 0.0014674874, 0.00744508, 0.011415428, 0.008664394, 0.0077569615, 0.007506847, 0.02971038, -8.9999998E15,
    0.82123715, 12.756191, 1.1000872, 0.9671487, 1.2557576, 6.3535967, 1.9879777, 6.0378857, 5.8721385, 0.29368687, 0.08297366, 1.2943926, 1.3520756, 9.051786, 2.0188982, 16.952885, 9.056293, 9.399705, 14.440703, -8.9999998E15,
    2.142261, 14.996106, 5.313879, 3.0252364, 9.933393, 16.23151, 11.753644, 11.43945, 8.575498, 0.2237048, 0.056117006, 5.0909204, 2.9520264, 3.7912745, 4.098896, 7.1546636, 5.000048, 4.010376, 12.19778, -8.9999998E15,
    3.098789, 19.561607, 14.097523, 13.047494, 14.250788, 12.508534, 14.091965, 8.301886, 5.8725004, 0.09821253, 0.036621276, 4.0736637, 2.3576517, 2.1588054, 3.0272002, 2.892411, 2.4637508, 2.223096, 6.7882595, -8.9999998E15,
    2.43078, 17.148699, 14.610028, 14.382902, 14.76154, 14.101113, 14.827712, 6.8873587, 4.3163486, 0.10815185, 0.024836391, 7.233815, 2.5374594, 0.9709879, 1.4043174, 0.60123014, 1.3285706, 1.032546, 2.658216, -8.9999998E15 ;
}
