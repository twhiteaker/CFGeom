netcdf nwm_bullcreek {
  dimensions:
    time = 1;
    station = 20;
  variables:
    int time(time);
      time:units = "seconds since 2016-05-26 06:00 UTC";
      time:long_name = "valid output time";

    int station_id(station);
      station_id:long_name = "Station id";

    double streamflow(station);
      streamflow:long_name = "River Flow";
      streamflow:units = "meter^3 / sec";

  // global attributes:
  :Conventions = "Unidata Observation Dataset v1.0";
  :cdm_datatype = "Station";
  :model_initialization_time = "2016-05-26_06:00:00";
  :station_dimension = "station";
  :missing_value = -8.9999998E15f;
  :stream_order_output = 1;
  :model_output_valid_time = "2016-05-27_00:00:00";
 data:

 time = 21600 ;

 station_id = 5781157, 5781193, 5781183, 5781189, 5781173, 5781133, 5781163, 
    5781131, 5781141, 5781171, 5781159, 5781129, 5781139, 5781149, 5781185, 
    5781187, 5781145, 5781781, 5781191, 5781811 ;

 streamflow = 0.252176284790039, 0.0201607346534729, 0.0346982032060623, 
    0.0607489943504334, 0.0835541933774948, 0.356544077396393, 
    0.105495147407055, 0.0702902525663376, 0.216611877083778, 
    0.0352071598172188, 0.0369682908058167, 0.101938299834728, 
    0.12274756282568, 0.375413328409195, 0.629893124103546, 
    0.717454493045807, 1.10981106758118, 1.15975689888, 1.37934672832489, 
    -1.99939995115805e-011 ;
}
