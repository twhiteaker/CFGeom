netcdf hucPolygons {
dimensions:
	maxStrlen64 = 64 ;
	station = 2 ;
	time = 25 ;
	char = 38 ;
	node = 2628 ;
variables:
	double lat(station) ;
		lat:units = "degrees_north" ;
		lat:missing_value = -999. ;
		lat:long_name = "latitude of the observation" ;
		lat:standard_name = "latitude" ;
    lat:nodes = "Y" ;
	double lon(station) ;
		lon:units = "degrees_east" ;
		lon:missing_value = -999. ;
		lon:long_name = "longitude of the observation" ;
		lon:standard_name = "longitude" ;
    lon:nodes = "X" ;
	double time(time) ;
		time:units = "days since 1970-01-01 00:00:00" ;
		time:missing_value = -999. ;
		time:long_name = "time of measurement" ;
		time:standard_name = "time" ;
	char station_name(station, maxStrlen64) ;
		station_name:units = "" ;
		station_name:missing_value = "" ;
		station_name:long_name = "Station Names" ;
		station_name:cf_role = "timeseries_id" ;
		station_name:standard_name = "station_id" ;
	int et(station, time) ;
		et:units = "mm" ;
		et:missing_value = -999 ;
		et:long_name = "Area Weighted Mean Actual Evapotranspiration" ;
		et:coordinates = "time lat lon" ;
		et:geometry = "geometry_container" ;
    et:grid_mapping = "crs" ;
	char TNMID(station, char) ;
		TNMID:units = "unknown" ;
	char METASOURCE(station, char) ;
		METASOURCE:units = "unknown" ;
	char SOURCEDATA(station, char) ;
		SOURCEDATA:units = "unknown" ;
	char SOURCEORIG(station, char) ;
		SOURCEORIG:units = "unknown" ;
	char SOURCEFEAT(station, char) ;
		SOURCEFEAT:units = "unknown" ;
	char LOADDATE(station, char) ;
		LOADDATE:units = "unknown" ;
	char GNIS_ID(station, char) ;
		GNIS_ID:units = "unknown" ;
	double AREAACRES(station) ;
		AREAACRES:units = "unknown" ;
		AREAACRES:_FillValue = NaN ;
		AREAACRES:geometry = "geometry_container" ;
    AREAACRES:grid_mapping = "crs" ;
	double AREASQKM(station) ;
		AREASQKM:units = "unknown" ;
		AREASQKM:_FillValue = NaN ;
		AREASQKM:geometry = "geometry_container" ;
    AREASQKM:grid_mapping = "crs" ;
	char STATES(station, char) ;
		STATES:units = "unknown" ;
	char HUC12(station, char) ;
		HUC12:units = "unknown" ;
	char NAME(station, char) ;
		NAME:units = "unknown" ;
	char HUTYPE(station, char) ;
		HUTYPE:units = "unknown" ;
	char HUMOD(station, char) ;
		HUMOD:units = "unknown" ;
	char TOHUC(station, char) ;
		TOHUC:units = "unknown" ;
	double NONCONTRIB(station) ;
		NONCONTRIB:units = "unknown" ;
		NONCONTRIB:_FillValue = NaN ;
		NONCONTRIB:geometry = "geometry_container" ;
    NONCONTRIB:grid_mapping = "crs" ;
	double NONCONTR_1(station) ;
		NONCONTR_1:units = "unknown" ;
		NONCONTR_1:_FillValue = NaN ;
		NONCONTR_1:geometry = "geometry_container" ;
    NONCONTR_1:grid_mapping = "crs" ;
	double SHAPE_Leng(station) ;
		SHAPE_Leng:units = "unknown" ;
		SHAPE_Leng:_FillValue = NaN ;
		SHAPE_Leng:geometry = "geometry_container" ;
    SHAPE_Leng:grid_mapping = "crs" ;
	double SHAPE_Area(station) ;
		SHAPE_Area:units = "unknown" ;
		SHAPE_Area:_FillValue = NaN ;
		SHAPE_Area:geometry = "geometry_container" ;
    SHAPE_Area:grid_mapping = "crs" ;
	double x(node) ;
		x:units = "degrees_east" ;
		x:standard_name = "longitude" ;
		x:axis = "X" ;
	double y(node) ;
		y:units = "degrees_north" ;
		y:standard_name = "latitude" ;
		y:axis = "Y" ;
	float geometry_container ;
		geometry_container:geometry_type = "polygon" ;
		geometry_container:node_count = "node_count" ;
		geometry_container:node_coordinates = "x y" ;
		geometry_container:coordinates = "lon lat" ;
		geometry_container:grid_mapping = "crs" ;
	int node_count(station) ;
		node_count:long_name = "count of coordinates in each instance geometry" ;
	float crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;
		crs:longitude_of_prime_meridian = 0. ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:featureType = "timeSeries" ;
		:cdm_data_type = "Station" ;
		:standard_name_vocabulary = "CF-1.7" ;
		:DODS.strlen = 12 ;
		:DODS.dimName = "name_strlen" ;
data:

 lat = 36.488959, 36.43594 ;

 lon = -80.399735, -80.365249 ;

 time = 10957, 10988, 11017, 11048, 11078, 11109, 11139, 11170, 11201, 11231, 
    11262, 11292, 11323, 11354, 11382, 11413, 11443, 11474, 11504, 11535, 
    11566, 11596, 11627, 11657, 11688 ;

 station_name =
  "030101030106",
  "030101030107" ;

 et =
  10, 19, 21, 36, 105, 110, 128, 121, 70, 25, 18, 9, 14, 17, 20, 54, 93, 127, 
    144, 125, 78, 29, 12, 9, 16,
  10, 20, 23, 37, 107, 114, 134, 118, 70, 27, 20, 8, 17, 20, 22, 61, 97, 133, 
    146, 123, 78, 30, 14, 11, 16 ;

 TNMID =
  "{94745C74-B81F-42C7-9397-09DE87E038D4}",
  "{D756B24D-1959-4938-8930-FC3D417BB708}" ;

 METASOURCE =
  "{2A42A390-4EEB-411B-928E-188529D9691D}",
  "NA" ;

 SOURCEDATA =
  "NA",
  "NA" ;

 SOURCEORIG =
  "NA",
  "NA" ;

 SOURCEFEAT =
  "NA",
  "NA" ;

 LOADDATE =
  "2013/01/18",
  "2013/01/18" ;

 GNIS_ID =
  "NA",
  "NA" ;

 AREAACRES = 28635, 8464 ;

 AREASQKM = 115.880118, 34.25262304 ;

 STATES =
  "NC",
  "NC" ;

 HUC12 =
  "030101030106",
  "030101030107" ;

 NAME =
  "Big Creek",
  "Double Creek" ;

 HUTYPE =
  "S",
  "S" ;

 HUMOD =
  "NM",
  "NM" ;

 TOHUC =
  "030101030109",
  "030101030109" ;

 NONCONTRIB = 0, 0 ;

 NONCONTR_1 = 0, 0 ;

 SHAPE_Leng = 0.668434563762557, 0.37395257288014 ;

 SHAPE_Area = 0.011654299957017, 0.003442696475335 ;

 x = -80.4339739845491, -80.4343932991317, -80.4346544887147, 
    -80.4349137376726, -80.4353912324635, -80.4358732980878, 
    -80.435980053296, -80.4362165491289, -80.4365028012118, 
    -80.4367297980864, -80.4368087387113, -80.436815930378, 
    -80.4368984897529, -80.4370954887109, -80.4373529845438, 
    -80.4373893657938, -80.43767073871, -80.4381968043342, -80.438516678292, 
    -80.4387451782916, -80.4388824887081, -80.4391676105827, 
    -80.4400202387063, -80.4404317355807, -80.4408374241218, 
    -80.4413196105793, -80.4416935480787, -80.4419592970366, 
    -80.442359109536, -80.4428711116186, -80.4433740543261, 
    -80.4436973605756, -80.4438244209921, -80.4444169886995, 
    -80.4453631095314, -80.445783924114, -80.4463383553632, -80.446711554321, 
    -80.4469626751539, -80.4472964866117, -80.4473213647367, 
    -80.4475647397363, -80.4483037959852, -80.4486649855679, 
    -80.4495267376499, -80.4501969230656, -80.4507785543147, 
    -80.4508628616062, -80.4508869251478, -80.4509108626478, 
    -80.4513558011888, -80.4518271084797, -80.4522162991041, 
    -80.4526293668118, -80.4530303678528, -80.4531574251443, 
    -80.4533050543107, -80.4534186751439, -80.4536043584769, 
    -80.4538729241015, -80.4541383605595, -80.4542094261843, 
    -80.454606050142, -80.4549781730581, -80.4553638001408, 
    -80.4556127376405, -80.4557491126403, -80.4557607397236, 
    -80.4557775459735, -80.4557720480569, -80.4558648001401, 
    -80.456141049098, -80.4565904251389, -80.4566482470138, 
    -80.4570347386799, -80.4573721793044, -80.4574908626375, 
    -80.4576341751373, -80.4578116740954, -80.4578943636786, 
    -80.4580389886784, -80.4582901740947, -80.4585354813859, 
    -80.4592995511764, -80.4600564220086, -80.4604343605496, 
    -80.4607394220075, -80.460823426174, -80.461493985548, -80.4619308001307, 
    -80.4624036157549, -80.4627583022127, -80.4631833001287, 
    -80.4635844865865, -80.4639494845025, -80.464277425127, 
    -80.4643256751269, -80.4648609251261, -80.4655586105417, 
    -80.4660756115825, -80.4665299907485, -80.4670716126227, 
    -80.4675847386636, -80.4680104272045, -80.4682276115792, 
    -80.4687131136618, -80.4691508636611, -80.4694471136607, 
    -80.469660989702, -80.4699575490765, -80.4702416167844, 
    -80.4705726199089, -80.470773487617, -80.4709627386583, 
    -80.4710581136582, -80.4710593615748, -80.4710724855332, 
    -80.4710732969915, -80.471168735533, -80.4714951771991, 
    -80.4720041094901, -80.4723223011562, -80.4723648646978, 
    -80.4728228667804, -80.4729362355303, -80.472897920947, -80.472879177197, 
    -80.4729537417802, -80.4731374886549, -80.4734004865712, 
    -80.4735657386543, -80.4735849271959, -80.4735795459459, 
    -80.4735617990709, -80.4736181740709, -80.4736669230291, 
    -80.473758304279, -80.4738204886539, -80.4741390511534, 
    -80.4743991115697, -80.4746359865693, -80.4749444240688, 
    -80.4751440511518, -80.4753477959432, -80.4757153615676, 
    -80.4761809834419, -80.47631292615, -80.4767044261494, -80.476753674066, 
    -80.47741611469, -80.4782070511471, -80.4788158605211, -80.4794751126034, 
    -80.4798550448945, -80.4801372980191, -80.4803958667687, 
    -80.4806666126016, -80.4809959865594, -80.4812897386423, 
    -80.4816352407251, -80.4817921782249, -80.4818009875998, 
    -80.4817044865583, -80.4816556761417, -80.4817130490583, 
    -80.4820286740578, -80.4822067396825, -80.4826666136402, 
    -80.4832216125976, -80.4837060490552, -80.4840721750963, 
    -80.4841896782211, -80.4841886678045, -80.4841981094711, 
    -80.4842150521794, -80.4842191146794, -80.4842404271794, 
    -80.484298050096, -80.4844386105124, -80.4848389907201, -80.485345860511, 
    -80.4856877990521, -80.4859474219684, -80.4862772355095, 
    -80.4864299261343, -80.4866063553007, -80.4868424230087, 
    -80.4875629896742, -80.48814142509, -80.4887549855057, -80.489398175088, 
    -80.4899517355038, -80.4902291125867, -80.4904676782114, 
    -80.4907861125859, -80.4910058615439, -80.4911259875853, 
    -80.4910873636271, -80.4909699282106, -80.4909117980023, 
    -80.4909525511273, -80.4911288021687, -80.4911517365437, 
    -80.4915137386264, -80.4921107386255, -80.4926535542497, 
    -80.4932434240404, -80.4934911761234, -80.4937508604979, 
    -80.4939048011227, -80.4940361157059, -80.4941440469557, 
    -80.4942086136222, -80.4944056740386, -80.4946791115382, 
    -80.4951308594542, -80.4954406136203, -80.4956068021617, 
    -80.4959501771612, -80.4965416073686, -80.4970881136177, 
    -80.4971331761177, -80.4975829907003, -80.4980337969496, 
    -80.4983546136158, -80.4990318021564, -80.4994114261142, 
    -80.4998616719468, -80.5006306729873, -80.5012569854863, 
    -80.5017531771522, -80.5019780511101, -80.5020731781934, 
    -80.5019680521519, -80.5018405500687, -80.5017492969439, 
    -80.5017676104855, -80.5020714865267, -80.5023565511096, 
    -80.5028672979838, -80.50317580215, -80.503580737566, -80.5040269250653, 
    -80.5045113000646, -80.5050311125638, -80.505503862563, 
    -80.5057524886043, -80.5059543021457, -80.5060262396456, 
    -80.5061225479787, -80.5062424219369, -80.5065042354781, 
    -80.5068133042276, -80.507240051102, -80.5077843604761, 
    -80.5084249896418, -80.5092271115156, -80.5097143594315, 
    -80.5101660427641, -80.5110419896378, -80.5118619271365, 
    -80.5119711083863, -80.5120334844279, -80.5120721750528, 
    -80.5121134198444, -80.5121559260944, -80.5121732313027, 
    -80.5122488010942, -80.5120513031779, -80.5120423615112, 
    -80.5121497990111, -80.512627050052, -80.5133919250508, 
    -80.5135919875505, -80.5138965521334, -80.5140106729665, 
    -80.5139779896332, -80.5137996750502, -80.5135918031755, 
    -80.5134356135924, -80.5128736104683, -80.5122348031776, 
    -80.5118976177615, -80.5115743635953, -80.5112328615125, 
    -80.5111636740126, -80.5107272375549, -80.5103056760972, 
    -80.5101513635975, -80.5098931094312, -80.5096554208899, 
    -80.5094906760985, -80.5092840510988, -80.5089258625577, 
    -80.5081043021423, -80.5077192333929, -80.5073766761018, 
    -80.507013486519, -80.5068538636026, -80.506816865686, -80.5069258656858, 
    -80.5065866125614, -80.5056560542295, -80.5050547365221, 
    -80.5045929250645, -80.5043470542315, -80.5038094886073, 
    -80.5032670511082, -80.5028602979838, -80.5022726761097, 
    -80.5019261125686, -80.5016097365274, -80.5015236115275, 
    -80.5011728011114, -80.5007208021538, -80.5001482959047, 
    -80.4999129250717, -80.4996357990305, -80.4989452969482, 
    -80.4988358636151, -80.4986748636153, -80.4986732354903, 
    -80.4986698604903, -80.4986208615321, -80.4984829250739, 
    -80.4979542375747, -80.4977702979917, -80.4972698625758, 
    -80.4970789865345, -80.4965797396602, -80.4964217334104, 
    -80.4962176729941, -80.4958268011197, -80.4956263615367, 
    -80.495198865704, -80.4947206782048, -80.4942671761222, 
    -80.4938506761228, -80.4935592375816, -80.4932159219571, 
    -80.4919727980007, -80.4912488605018, -80.4904104209198, 
    -80.4897155532125, -80.4891463605051, -80.4891179271718, 
    -80.4888332375889, -80.488516863631, -80.4881552396733, 
    -80.4876881719657, -80.4874278657161, -80.4872361750914, 
    -80.4868444855086, -80.4866184928007, -80.4864075480094, 
    -80.4861061761348, -80.4855788698856, -80.485126861553, 
    -80.4846598000954, -80.4841927375961, -80.4836654271803, 
    -80.4832254813476, -80.4831229855145, -80.4827312990567, 
    -80.4824751719738, -80.4824241084322, -80.4823094250991, 
    -80.4820637344744, -80.4819477980163, -80.4815561751002, 
    -80.480802738643, -80.4802603584355, -80.4799288657277, 
    -80.4797782355196, -80.479778240728, -80.4797933001029, 
    -80.4797330501031, -80.4795974251032, -80.4792508626038, 
    -80.4789194219793, -80.4784824886466, -80.4781058001056, 
    -80.4779250490642, -80.4776839907312, -80.4775494219815, 
    -80.4773374271901, -80.4772601761485, -80.4769411740657, 
    -80.4768747334408, -80.4767322407327, -80.475902734484, 
    -80.4751353021935, -80.4746441782359, -80.4739686115703, 
    -80.4739661042786, -80.4736009271959, -80.4732844865714, 
    -80.4731489271966, -80.4730434188634, -80.4728928001136, 
    -80.4727708636555, -80.4722948532396, -80.4718792376152, 
    -80.4717506730321, -80.4717143011571, -80.4712089261579, 
    -80.4708256136585, -80.4706041740756, -80.4704218636592, 
    -80.4702410490761, -80.4699547376182, -80.4696685542853, 
    -80.4694877397023, -80.4692617376193, -80.469020674078, 
    -80.4687042324118, -80.4683878626207, -80.4678304209548, 
    -80.4676306147052, -80.467272929289, -80.4669113636646, -80.46662504804, 
    -80.466431552207, -80.466203175124, -80.4659169199162, -80.4656352438749, 
    -80.4654799865835, -80.4650279876258, -80.4645910501266, 
    -80.4644554865851, -80.46448561471, -80.4645662376266, -80.4646513605431, 
    -80.4648170542928, -80.4648623074178, -80.4648019897095, 
    -80.4645759865849, -80.4642445511687, -80.4637323053362, 
    -80.4636964220029, -80.4632351188786, -80.4628433605459, 
    -80.4625721792963, -80.4623160511717, -80.4620146772139, 
    -80.4613066105483, -80.4610673647153, -80.4609569292989, 
    -80.4608582928407, -80.4608002970074, -80.4605840501328, 
    -80.4598148615923, -80.4591829834683, -80.4587498043023, 
    -80.458495050136, -80.4580816813867, -80.4577721126371, 
    -80.4575399251375, -80.4573289865962, -80.4571783022214, 
    -80.4570426772216, -80.4569673626384, -80.4568318053469, 
    -80.4566811115972, -80.4564701730558, -80.4561085532647, 
    -80.4556867365987, -80.4553853626408, -80.455249803266, 
    -80.4552497949327, -80.4553853626408, -80.4553979907658, 
    -80.4554154865991, -80.4553251168076, -80.4551744230578, 
    -80.4549032428499, -80.4547073636836, -80.4545567313921, 
    -80.4544964209755, -80.4544964209755, -80.4544964188922, 
    -80.4543909876423, -80.454180052226, -80.4538786741015, 
    -80.4538739897265, -80.4535321761854, -80.4531706084776, 
    -80.4526733636867, -80.4521008595209, -80.4516488626466, 
    -80.4514981709802, -80.4514529866053, -80.4514981751469, 
    -80.4516639241049, -80.4517396720215, -80.4517995522297, 
    -80.4517995543131, -80.4517392386882, -80.4515433657718, 
    -80.451181801189, -80.4506695491065, -80.4503229876487, 
    -80.4501421782739, -80.4499764866076, -80.4497956709828, 
    -80.4496751126497, -80.449675114733, -80.4496751105664, 
    -80.4495997980665, -80.4494189876501, -80.4491176772339, 
    -80.4488012959844, -80.4483341772351, -80.4480821751521, 
    -80.4478671116108, -80.4475356136947, -80.4472795501534, 
    -80.446917925154, -80.446722113696, -80.4465714261962, -80.4464809886963, 
    -80.4465111751546, -80.4466768647377, -80.4470083657789, 
    -80.447108111612, -80.4473548605699, -80.4478822418191, 
    -80.4482287355686, -80.44839448661, -80.4483944886933, -80.4482437980686, 
    -80.4481512991104, -80.447927426194, -80.4476562366112, 
    -80.4474001116116, -80.4473601116116, -80.4472481772368, 
    -80.4469136761957, -80.4467006751543, -80.4463950480715, 
    -80.4463642386965, -80.4463303605716, -80.4461797376551, 
    -80.4459235480722, -80.4456523616143, -80.4453811720314, 
    -80.4450948605735, -80.4448237355739, -80.444541424116, 
    -80.4444621105744, -80.4440854209917, -80.4437690501588, 
    -80.4433773012011, -80.4429704939101, -80.4428348616186, 
    -80.4427143647438, -80.4426511137023, -80.4424883605775, 
    -80.4422171730779, -80.4419610480783, -80.4419309230784, 
    -80.4419139262034, -80.4418856782868, -80.4418856699534, 
    -80.4417952980786, -80.4415994241206, -80.4412981105793, 
    -80.4410118626631, -80.440695427247, -80.4402735470393, 
    -80.4398667959982, -80.4397462376651, -80.4397161137068, 
    -80.4398969241232, -80.4401379897478, -80.4405447355805, 
    -80.4407948626635, -80.4409515522466, -80.4413734220376, 
    -80.4415693001623, -80.4417953001619, -80.4418555491201, 
    -80.4418404866202, -80.4417501084953, -80.4417055512037, 
    -80.4416747355788, -80.441719984537, -80.4418404876619, 
    -80.4420295480782, -80.4422171741196, -80.4426088605773, 
    -80.4429554251601, -80.4432115512014, -80.4434224887011, 
    -80.4434375522427, -80.4433170501596, -80.4431211699516, 
    -80.442849985577, -80.4426842366189, -80.4425335564108, -80.442413047036, 
    -80.4421417282864, -80.4417651762037, -80.4415090470374, 
    -80.4413975491209, -80.441087175163, -80.4406201147471, 
    -80.4403171720392, -80.4402983022476, -80.4401684209978, 
    -80.4401032980812, -80.4399119876649, -80.4397914262067, 
    -80.4397311751652, -80.4397311751652, -80.4395955501653, 
    -80.4393846126657, -80.4392038637076, -80.4391887980826, 
    -80.4393092991241, -80.4394736730822, -80.4395202376655, 
    -80.4397462376651, -80.4398818626649, -80.4398667991233, 
    -80.4395653637071, -80.4392189272493, -80.4388723626665, 
    -80.4385258605836, -80.4381039887093, -80.4376067980851, 
    -80.4372903626689, -80.4368383605863, -80.4365370564201, 
    -80.4362959876705, -80.4360785460041, -80.4360399262125, 
    -80.4357837355879, -80.43554267413, -80.4352262355888, -80.4348043668394, 
    -80.4342318605903, -80.4336291157996, -80.4330717376754, 
    -80.4325896126762, -80.4320321116354, -80.4316554845527, 
    -80.431203485595, -80.4306911762208, -80.4300433637218, 
    -80.4299822991386, -80.4294256730978, -80.4290037408068, 
    -80.428878234557, -80.4285216105992, -80.4279189314335, 
    -80.4273614866427, -80.4270601699765, -80.4266985460187, 
    -80.4258849262283, -80.4250562991463, -80.4246946741468, 
    -80.4243632366473, -80.4242902991474, -80.4242794866474, 
    -80.423479738732, -80.4217203626931, -80.4210482366524, 
    -80.4208697376944, -80.4201158564456, -80.4196963022795, 
    -80.4196514897797, -80.4196129251964, -80.41937086478, -80.4189723595724, 
    -80.4186159887396, -80.4180586126988, -80.4173447397832, 
    -80.4164515502013, -80.4157956814523, -80.4149439241619, 
    -80.4134414252059, -80.4127701147903, -80.4123173627077, 
    -80.4120230481248, -80.4118077356251, -80.4115515512505, 
    -80.4112712387509, -80.4112543647927, -80.4109568054181, 
    -80.4105616137521, -80.4101871731277, -80.4100707991695, 
    -80.4097554845866, -80.4091728606292, -80.4087787377132, 
    -80.4085388033386, -80.4083331731305, -80.4080761762559, 
    -80.407789986673, -80.4073601752154, -80.4063725502169, 
    -80.4061852387588, -80.4057195523013, -80.404768738761, 
    -80.4040361731372, -80.4031067398053, -80.4025720543895, 
    -80.4018990502238, -80.401365611683, -80.4009024273087, 
    -80.4007590502256, -80.4005534221009, -80.4003477991846, 
    -80.4001764241848, -80.4000050533518, -80.3998508710604, 
    -80.3997436127272, -80.3996424877274, -80.3994022991861, 
    -80.3993873668944, -80.3986858054372, -80.3976923616887, 
    -80.3965413627321, -80.3957283012751, -80.3948172346098, 
    -80.3944759273187, -80.3944406148187, -80.3939654231528, 
    -80.3936612377366, -80.3935619252368, -80.3934076741954, 
    -80.3933221189872, -80.3930992408625, -80.392585173155, 
    -80.3921568012806, -80.3917454887813, -80.391282863782, 
    -80.3910429231574, -80.3909743606575, -80.3909059273242, 
    -80.3908591137827, -80.3907858648244, -80.3906830471163, 
    -80.3903917367001, -80.3896891710762, -80.3892359856602, 
    -80.3889711700356, -80.3887328012859, -80.388699054411, -80.388690985661, 
    -80.3885306752446, -80.3877361117042, -80.3875981137877, 
    -80.3875814221211, -80.3869474210804, -80.3866217992059, 
    -80.3865018627478, -80.3863990492063, -80.3864161762896, 
    -80.3866903669141, -80.3867611752473, -80.386528674206, 
    -80.3862584283732, -80.3859488606653, -80.3856604210824, 
    -80.3853712919162, -80.3851054867083, -80.3848904887919, 
    -80.3845902356674, -80.3838107398353, -80.3834190492109, 
    -80.3831324856696, -80.382515922129, -80.3823408627542, 
    -80.3820232377547, -80.3815093617138, -80.3814712981722, 
    -80.3807166158817, -80.3802219231741, -80.3800879262994, 
    -80.3796303023418, -80.3792190513007, -80.3787735450514, 
    -80.3784136752603, -80.3783482367188, -80.3782769200522, 
    -80.3781534263024, -80.378150989844, -80.3782866763022, 
    -80.3783237388021, -80.3780851773441, -80.3778438638029, 
    -80.3773857950536, -80.3770274221375, -80.3768299273461, 
    -80.3768341106794, -80.3767970502628, -80.376717800263, 
    -80.3763633606802, -80.3757504856811, -80.3751171763071, 
    -80.3748995585991, -80.3746818617244, -80.3740306096421, 
    -80.3738089888091, -80.3737359877676, -80.3735016763096, 
    -80.3732874242266, -80.3729344252688, -80.3722266721449, 
    -80.3717537981873, -80.3713413586046, -80.3710772981884, 
    -80.3707024242306, -80.3704282971477, -80.3701712992314, 
    -80.369571484649, -80.3691259283997, -80.3685947356922, 
    -80.3681694211095, -80.3679606836099, -80.3677207992353, 
    -80.3674466159023, -80.367001050278, -80.3667152367368, -80.366589802362, 
    -80.3661956690293, -80.3658529273631, -80.3653731752805, 
    -80.3647733627815, -80.3644649252819, -80.3643981773654, 
    -80.3643054888238, -80.3642908034072, -80.3642421846573, 
    -80.3641790534074, -80.3641517992407, -80.3641393648658, 
    -80.3641222377825, -80.3641164221575, -80.3640867388242, 
    -80.3638474898663, -80.3634706117418, -80.3632118638255, 
    -80.362927363826, -80.3628399252845, -80.3627389232013, 
    -80.3620842377857, -80.3615892357031, -80.3613126742452, 
    -80.3608801086208, -80.3605683586213, -80.3603284242467, 
    -80.3600687357055, -80.3597583659143, -80.3596464200811, 
    -80.3594662357063, -80.3593249263316, -80.3591634252902, 
    -80.3590209200821, -80.3588019252907, -80.3585625492494, 
    -80.3584027971664, -80.3581251107084, -80.3573741763346, 
    -80.3569391773769, -80.3563654273779, -80.3559301752952, 
    -80.3554562377959, -80.3553274867544, -80.3552429315463, 
    -80.3552201815463, -80.355197604463, -80.3550927971715, 
    -80.3549853596717, -80.3548693617552, -80.3546529909222, 
    -80.354317608631, -80.353903235715, -80.353509365924, -80.3531566107162, 
    -80.3530355482164, -80.3525216784255, -80.3521701763427, 
    -80.3519876096763, -80.3515339878021, -80.3514142325939, 
    -80.351121111761, -80.3504314232204, -80.3500224253044, 
    -80.3499584211378, -80.3498942378046, -80.349427301347, 
    -80.3488356732229, -80.3481841711405, -80.3478980503077, 
    -80.3471756773921, -80.3464452336433, -80.3458733721858, 
    -80.3453770513532, -80.34532041802, -80.3444324930214, -80.3434838596895, 
    -80.3430091773986, -80.3426319836492, -80.3421557357332, 
    -80.3416210524007, -80.340570175319, -80.3396368044872, 
    -80.3390010513631, -80.3386230524054, -80.3385746680304, 
    -80.3383631774058, -80.3381239242811, -80.3377270503235, 
    -80.3374427961572, -80.3371325544911, -80.3367162399084, 
    -80.3364967992837, -80.3364158024089, -80.3363932982422, 
    -80.3362747409507, -80.3362524242841, -80.3361269899092, 
    -80.3359932899095, -80.3356542357433, -80.3352970513689, -80.33460398887, 
    -80.334108234704, -80.3338917992878, -80.3332196753304, 
    -80.3329440534559, -80.3327874867895, -80.3326813628313, 
    -80.3325920544981, -80.3317837357494, -80.3304908628347, 
    -80.3304648617931, -80.3298548545023, -80.329046109712, 
    -80.3289436732538, -80.3286127367959, -80.3281596784633, 
    -80.3278239232555, -80.3273427347146, -80.3271769242982, 
    -80.3267142399239, -80.326200173258, -80.3256861732588, 
    -80.3252405503428, -80.3250563024264, -80.3248766763851, 
    -80.3245209836773, -80.3245071743023, -80.3241844857611, 
    -80.3239989243031, -80.3239039253449, -80.3238182357617, 
    -80.3235612305538, -80.3233556107624, -80.3232022961793, 
    -80.3230299868046, -80.3227215493051, -80.3226016138886, 
    -80.3224816722221, -80.3222759878474, -80.3220499847228, 
    -80.3220361055562, -80.3219901690979, -80.3216419888901, 
    -80.3212478607657, -80.3207884243081, -80.3205981732667, 
    -80.3204810503502, -80.3201381128508, -80.3200882368092, 
    -80.3196743586848, -80.319556796185, -80.319360425352, -80.3186493618114, 
    -80.3180450513957, -80.3174607972299, -80.3171009232722, 
    -80.3167582388976, -80.3164154868149, -80.3162784222317, 
    -80.3163297972317, -80.3163812378566, -80.3162716732734, 
    -80.3162378607735, -80.315925854524, -80.3155094899413, 
    -80.3149219264005, -80.3149215503589, -80.3144874847345, 
    -80.313973173277, -80.3134186711945, -80.3130238014035, 
    -80.3128468628621, -80.3126819222373, -80.3125381107792, 
    -80.3126503597374, -80.3127207972373, -80.3129882993202, 
    -80.3130911139034, -80.3130911097367, -80.3131596753616, 
    -80.313279607653, -80.3133824274446, -80.3133824222363, 
    -80.3133138618197, -80.3131596743199, -80.3129539857786, 
    -80.3125770514042, -80.3122111764047, -80.312026926405, 
    -80.3110422357815, -80.310330240991, -80.3096986764086, 
    -80.3090403014097, -80.3084620493272, -80.3080287420363, 
    -80.3070466118294, -80.3063624941221, -80.3056871732899, 
    -80.3053653628737, -80.3050006732909, -80.3046407337081, 
    -80.3035253003765, -80.3028341139193, -80.3022611118369, 
    -80.3020554795455, -80.3019698014206, -80.3018498618375, 
    -80.3018111732958, -80.3015756712129, -80.3012329857968, 
    -80.3009073618389, -80.3005818045478, -80.3005132337145, 
    -80.3005475503812, -80.3005646764228, -80.3004447347563, 
    -80.3001536128818, -80.3001362399651, -80.299810670174, 
    -80.2994654899662, -80.2991554243417, -80.2987676149673, 
    -80.2983724858012, -80.2981543628849, -80.2980651774683, 
    -80.2981304858016, -80.2980182389268, -80.2978132941354, 
    -80.2970522951783, -80.2964995493458, -80.2956722368471, 
    -80.2948459805983, -80.2944820503906, -80.2935918681003, 
    -80.2931314910177, -80.2925267983103, -80.2918132410197, 
    -80.2912517983123, -80.2906428608132, -80.2900254253975, 
    -80.2889847399824, -80.2886264858163, -80.2885164243582, 
    -80.2884569274833, -80.2884484878999, -80.2880364243589, 
    -80.2876406045679, -80.2871462399853, -80.2868204264441, 
    -80.2864193014448, -80.2860957399869, -80.2859776201955, 
    -80.2857696764458, -80.2853430524881, -80.284747111864, 
    -80.2847071191558, -80.2847057618641, -80.2846275858225, 
    -80.2846992191558, -80.284948357697, -80.2853608629047, -80.285816241029, 
    -80.2861412399869, -80.2863994212365, -80.2867300483193, 
    -80.2868254295691, -80.2871171733187, -80.2876049233179, 
    -80.2880544879006, -80.2885446128998, -80.2887789233161, 
    -80.2889347389408, -80.2894058014401, -80.2898186108145, 
    -80.2899946733142, -80.290110235814, -80.2903644253969, 
    -80.2908744899795, -80.2912671128956, -80.2914028628954, 
    -80.2914210462287, -80.2914569878953, -80.2915736118534, 
    -80.2917902368531, -80.2923037983106, -80.2926596118517, 
    -80.2928172378932, -80.2931119920594, -80.2937039858085, 
    -80.2940577337246, -80.2941733628911, -80.294208422266, 
    -80.2942104264326, -80.2944658003906, -80.2942459243493, 
    -80.294184734766, -80.2943012358076, -80.294438555599, -80.2945670503905, 
    -80.2953552993475, -80.2959036743467, -80.2960578628881, 
    -80.2961435576797, -80.2962978649711, -80.2963662983043, 
    -80.2964862993458, -80.2964737972625, -80.2964348639292, 
    -80.2963834847626, -80.2964519910125, -80.2965034264291, 
    -80.2964519858042, -80.2964519889292, -80.2964519868459, 
    -80.2966233639289, -80.2969317920534, -80.2970346170533, 
    -80.2969661149701, -80.2967090493455, -80.2964177347626, 
    -80.2961264170547, -80.2957245514303, -80.2955952993472, 
    -80.2951838649728, -80.2949440514315, -80.2947555493485, 
    -80.2948069285151, -80.2949440514315, -80.2951496764312, 
    -80.2952696118477, -80.2952524868477, -80.2951496722645, 
    -80.2950982389313, -80.2950126097647, -80.2949611712232, 
    -80.2949783014315, -80.2951496774729, -80.2954067399725, 
    -80.2958008639302, -80.2962670503878, -80.2964863003875, 
    -80.2968804253869, -80.2971031712198, -80.2973773639278, 
    -80.2976344264274, -80.2977747368438, -80.2980799180933, 
    -80.2984055535095, -80.2988339285088, -80.299347984758, -80.299793548299, 
    -80.2999447316321, -80.30130455038, -80.3017825493376, -80.3020041076706, 
    -80.302141174337, -80.3021411764204, -80.3021411816287, 
    -80.3021411722537, -80.3023125472535, -80.3026552399612, 
    -80.3027066660028, -80.3026381149613, -80.3026381128779, 
    -80.3026552357945, -80.3027580482944, -80.3029808618357, 
    -80.3033749826685, -80.3037176764179, -80.3038469805844, 
    -80.3042317972505, -80.3044888014167, -80.3046772982914, 
    -80.3048315545412, -80.3048829222494, -80.3050371743325, 
    -80.3051057430824, -80.3050543024575, -80.3050001128743, 
    -80.3049515534993, -80.3048315503745, -80.3049515503743, 
    -80.3051913576656, -80.3054141753736, -80.3059111139145, 
    -80.3059869232894, -80.3064080420388, -80.3064252337054, 
    -80.3064937347469, -80.3065279847469, -80.3067336191216, 
    -80.3072477368291, -80.3076438639118, -80.307933177453, 
    -80.3082587326609, -80.308618608702, -80.3089270534932, 
    -80.3091841128677, -80.3094068597424, -80.3094833618256, 
    -80.3096639264087, -80.309886674325, -80.3100237378665, 
    -80.3101951159912, -80.3103835482826, -80.3107777378653, 
    -80.3111376180731, -80.3115488597391, -80.3121486097381, 
    -80.3125427378625, -80.3128683618204, -80.31313529932, -80.3140539264019, 
    -80.3150949868169, -80.3157147388993, -80.3160505493154, 
    -80.3160559899404, -80.3161859243152, -80.3161043013987, 
    -80.3158642347324, -80.3154658055664, -80.3153845441082, 
    -80.3154802368163, -80.3155073034829, -80.3155073034829, 
    -80.315455865983, -80.3153530503582, -80.3151988586918, 
    -80.3151816774418, -80.3153016753583, -80.3155586753579, 
    -80.3158499857741, -80.3160899295237, -80.3161934253569, 
    -80.3163641159816, -80.3164840503565, -80.3165011701481, 
    -80.3163812399399, -80.3162557326485, -80.3161242399403, 
    -80.3158671034824, -80.3158157388991, -80.3157643013992, 
    -80.3157814888992, -80.3159699232739, -80.3162955503567, 
    -80.3165868649396, -80.3168953003558, -80.317181238897, 
    -80.3176249201463, -80.3177412347295, -80.3176199847297, 
    -80.3177784284794, -80.318472863895, -80.3188414211861, 
    -80.3190776066024, -80.3190948638941, -80.3189746118109, 
    -80.3187561138946, -80.3183990524368, -80.318261236812, 
    -80.3176468013963, -80.3172685513969, -80.3170872368138, 
    -80.317004739939, -80.3170613003555, -80.3169597420223, 
    -80.3167593638977, -80.3166375451478, -80.3166749878561, 
    -80.3168706159808, -80.316987052439, -80.316965043064, -80.3170222972306, 
    -80.3174134857717, -80.3178841763959, -80.3183074941036, 
    -80.318510863895, -80.319081551394, -80.3192969836854, -80.3194133024352, 
    -80.3194094295185, -80.3192772357688, -80.3190887357691, 
    -80.3190030472275, -80.3190544263941, -80.3192943649354, 
    -80.3200140493093, -80.3202367993089, -80.3203567972254, 
    -80.3204424857669, -80.3206823649332, -80.3211964274324, 
    -80.3216248597234, -80.3220703638895, -80.3224644826388, 
    -80.3228322378466, -80.3228757993048, -80.3232528003459, 
    -80.3235441107622, -80.3237154253452, -80.3238525482616, 
    -80.3239382409699, -80.3241007357612, -80.3245248024273, 
    -80.3250004826349, -80.325338236801, -80.325755362842, -80.326628555549, 
    -80.3274853597143, -80.3278109878389, -80.3280337357552, 
    -80.3282564878381, -80.3285306722127, -80.3286406732542, 
    -80.3288049242957, -80.3289419263788, -80.329010487837, 
    -80.3290104857537, -80.3288733597122, -80.3287864878373, 
    -80.328753426379, -80.3288733586705, -80.3289108628371, -80.32921611492, 
    -80.3296959263776, -80.3297301763776, -80.3297301763776, 
    -80.3296444857527, -80.3294731742946, -80.3292124284617, 
    -80.3291646795034, -80.328753426379, -80.328582049296, -80.3284449867962, 
    -80.3283936138796, -80.3284501690878, -80.3284324826295, 
    -80.3289077367955, -80.3292936117949, -80.3296582357527, 
    -80.3297109222109, -80.3299015565856, -80.3305356128346, 
    -80.3308782930424, -80.3310648628338, -80.3312724284585, 
    -80.3316298607496, -80.3316836763745, -80.3320435472073, 
    -80.3325233024149, -80.3330203013724, -80.3333972972052, 
    -80.3336373076215, -80.3337228628297, -80.3336200503298, 
    -80.3335686732466, -80.3336886128297, -80.3339970513709, 
    -80.3347168003281, -80.3349224211611, -80.3351452347025, 
    -80.3354022367854, -80.3354560451186, -80.3357106763683, 
    -80.3358991753263, -80.3361219253259, -80.3366784284501, 
    -80.3367731117833, -80.3374242982406, -80.3381610471978, 
    -80.3390179253215, -80.3399604242783, -80.3404830544858, 
    -80.3411428034432, -80.3413827336511, -80.3415198003175, 
    -80.341673988859, -80.3418796076087, -80.3421024232333, 
    -80.3423938023996, -80.3428049888573, -80.3431106148984, 
    -80.343387614898, -80.3438331742723, -80.3443129878132, 
    -80.3445186086462, -80.3447927357291, -80.3449469878122, 
    -80.3449998023955, -80.3450155492705, -80.3452554242701, 
    -80.3454468044781, -80.3455057961447, -80.3457214138527, 
    -80.3462001784353, -80.3471809846838, -80.3473542305168, 
    -80.3486577378065, -80.3489764888477, -80.3494372367636, 
    -80.3496765523882, -80.349830733638, -80.3499334857212, 
    -80.3499334898879, -80.3497279221799, -80.3496765513466, 
    -80.3496694857216, -80.3496594221799, -80.3496765471799, 
    -80.3498821721796, -80.3503449273872, -80.3507328013449, 
    -80.3510816711361, -80.3512530492608, -80.3514757971771, -80.35175004926, 
    -80.3521269836344, -80.3526581742586, -80.353292235716, 
    -80.3539091117566, -80.3542347357145, -80.3544746107141, 
    -80.3546631107138, -80.3550229888383, -80.3554513638376, 
    -80.3563081763363, -80.3570450502935, -80.3574563013345, 
    -80.3578161742506, -80.3580731784169, -80.3582788013332, 
    -80.3586557992493, -80.3589814284155, -80.359289859665, 
    -80.3593866169565, -80.3596154242478, -80.3597696752892, 
    -80.3600095471639, -80.3604037388299, -80.3610377367456, 
    -80.3616889263279, -80.3620144232024, -80.3623057971603, 
    -80.3624428638267, -80.3626484815348, -80.362905548201, 
    -80.3632996732004, -80.3636595471582, -80.3644306148653, 
    -80.3652267356974, -80.365287480489, -80.3658015502799, 
    -80.3661785471543, -80.3666628627785, -80.3671052356945, 
    -80.3677268023602, -80.3679853638181, -80.3684404856925, 
    -80.3690231179832, -80.3695714898574, -80.3699313638151, 
    -80.3700980544399, -80.3702226742313, -80.3704282971477, 
    -80.370668110689, -80.370890928397, -80.3713706763129, -80.3717821138123, 
    -80.3722446721449, -80.3728272981857, -80.3732900502683, 
    -80.3737012388093, -80.3741467961003, -80.3743866752666, 
    -80.3745338033913, -80.3746951763077, -80.374969296099, 
    -80.3752778002652, -80.375808985681, -80.3762257356804, 
    -80.3764919283883, -80.3768835450543, -80.3772581106788, 
    -80.3777119867197, -80.3783048627604, -80.3792948658839, 
    -80.3800879940077, -80.3806436742152, -80.3810726085895, 
    -80.3819436096298, -80.3821879231711, -80.3823202377542, 
    -80.3831426148363, -80.3833662356693, -80.3834924877524, 
    -80.3836424867105, -80.3848916721253, -80.3853883033745, 
    -80.3854058585828, -80.3855331762909, -80.3855906085825, 
    -80.3856274314991, -80.3857701804572, -80.385902236707, 
    -80.3860796106651, -80.38616173879, -80.3863184210813, -80.3868274856639, 
    -80.387392926288, -80.3877871742041, -80.3880955512869, 
    -80.3882668669117, -80.388506799203, -80.3887809887859, 
    -80.3890037387855, -80.3891751148269, -80.3893292992017, 
    -80.389530550243, -80.389534990868, -80.3895612356596, -80.389757736701, 
    -80.3901347398254, -80.3905974252414, -80.3908715502409, 
    -80.3911114887823, -80.391265673157, -80.3913684877402, 
    -80.3914884887816, -80.3917219856563, -80.3917724856562, 
    -80.3921895512806, -80.3927034252381, -80.3937653023198, 
    -80.3946138596102, -80.394692925235, -80.3948128606515, 
    -80.3950184919012, -80.3952926752341, -80.3956867971085, 
    -80.3960432439829, -80.3960449856496, -80.3965366148155, 
    -80.3967849866901, -80.3972728637727, -80.3982447346045, 
    -80.3987057991872, -80.399250365853, -80.3995779231441, 
    -80.3999256752269, -80.4003754231429, -80.4010968596001, 
    -80.4012618606415, -80.4015197418911, -80.4018726137655, 
    -80.4022032970984, -80.402450737723, -80.4037711148043, 
    -80.4054344866767, -80.406339553342, -80.4070107429242, 
    -80.4075330512568, -80.4079344210478, -80.4081234835475, 
    -80.408277606464, -80.4083967377138, -80.4084934252136, 
    -80.4086129210468, -80.4087154877133, -80.4087671116715, 
    -80.4091669283376, -80.4097270512534, -80.4102497377109, 
    -80.4108734877099, -80.4108823627099, -80.4114132981258, 
    -80.4119604845832, -80.4126172397906, -80.4130894887481, 
    -80.413407487706, -80.4134158022893, -80.4135591720807, 
    -80.4136038606223, -80.4135649908308, -80.4134787387475, 
    -80.4134312991643, -80.413381918956, -80.4131898002063, 
    -80.4131039262481, -80.4130778627065, -80.413146801248, 
    -80.4132866095812, -80.4133819856227, -80.4135147387475, 
    -80.4137127377055, -80.4143452377045, -80.4151875502032, 
    -80.4156958606191, -80.4159442335354, -80.4161813533267, 
    -80.416454988743, -80.4167991127007, -80.4172136147834, 
    -80.4173307991582, -80.4177692376992, -80.4181119251987, 
    -80.4185129293647, -80.4188069887393, -80.4191012345722, 
    -80.4195618043631, -80.4201406158205, -80.4204000470701, 
    -80.4207073001946, -80.4211801751939, -80.4215977397766, 
    -80.4218871762345, -80.4222644866506, -80.4226898022749, 
    -80.4233559908155, -80.4242624856058, -80.4255402345622, 
    -80.4258239866451, -80.4259532949782, -80.4259398637282, 
    -80.4259254856032, -80.4259462970615, -80.4260628033114, 
    -80.4263447428942, -80.4268276106018, -80.4270432387265, 
    -80.4280117991416, -80.4290663001817, -80.4296201147641, 
    -80.4300441158052, -80.4303146126798, -80.4305134262211, 
    -80.4305571147627, -80.4306398647626, -80.4307438022624, 
    -80.4308960522622, -80.4311672366367, -80.4315454230945, 
    -80.4317531116358, -80.431864238719, -80.432097928302, -80.4324551095514, 
    -80.4328955480924, -80.4331532376754, -80.433557299133, 
    -80.4339739845491, -80.2970522951783, -80.2978132941354, 
    -80.2980182389268, -80.2981304858016, -80.2980651774683, 
    -80.2981543628849, -80.2983724858012, -80.2987676149673, 
    -80.2991554243417, -80.2994654899662, -80.299810670174, 
    -80.3001362399651, -80.3001536128818, -80.3004447347563, 
    -80.3005646764228, -80.3005475503812, -80.3005132337145, 
    -80.3005818045478, -80.3009073618389, -80.3012329857968, 
    -80.3015756712129, -80.3018111732958, -80.3018498618375, 
    -80.3019698014206, -80.3020554795455, -80.3022611118369, 
    -80.3028341139193, -80.3035253003765, -80.3046407337081, 
    -80.3050006732909, -80.3053653628737, -80.3056871732899, 
    -80.3063624941221, -80.3070466118294, -80.3080287420363, 
    -80.3084620493272, -80.3090403014097, -80.3096986764086, 
    -80.310330240991, -80.3110422357815, -80.312026926405, -80.3122111764047, 
    -80.3125770514042, -80.3129539857786, -80.3131596743199, 
    -80.3133138618197, -80.3133824222363, -80.3133824274446, 
    -80.313279607653, -80.3131596753616, -80.3130911097367, 
    -80.3130911139034, -80.3129882993202, -80.3127207972373, 
    -80.3126503597374, -80.3125381107792, -80.3126819222373, 
    -80.3128468628621, -80.3130238014035, -80.3134186711945, 
    -80.313973173277, -80.3144874847345, -80.3149215503589, 
    -80.3149219264005, -80.3155094899413, -80.315925854524, 
    -80.3162378607735, -80.3162716732734, -80.3163812378566, 
    -80.3163297972317, -80.3162784222317, -80.3164154868149, 
    -80.3167582388976, -80.3171009232722, -80.3174607972299, 
    -80.3180450513957, -80.3186493618114, -80.319360425352, -80.319556796185, 
    -80.3196743586848, -80.3200882368092, -80.3201381128508, 
    -80.3204810503502, -80.3205981732667, -80.3207884243081, 
    -80.3212478607657, -80.3216419888901, -80.3219901690979, 
    -80.3220361055562, -80.3220499847228, -80.3222759878474, 
    -80.3224816722221, -80.3226016138886, -80.3227215493051, 
    -80.3230299868046, -80.3232022961793, -80.3233556107624, 
    -80.3235612305538, -80.3238182357617, -80.3239039253449, 
    -80.3239989243031, -80.3241844857611, -80.3245071743023, 
    -80.3245209836773, -80.3248766763851, -80.3250563024264, 
    -80.3252405503428, -80.3256861732588, -80.326200173258, 
    -80.3267142399239, -80.3271769242982, -80.3273427347146, 
    -80.3278239232555, -80.3281596784633, -80.3286127367959, 
    -80.3289436732538, -80.329046109712, -80.3298548545023, 
    -80.3304648617931, -80.3304908628347, -80.3317837357494, 
    -80.3325920544981, -80.3326813628313, -80.3327874867895, 
    -80.3329440534559, -80.3332196753304, -80.3338917992878, 
    -80.334108234704, -80.33460398887, -80.3352970513689, -80.3356542357433, 
    -80.3359932899095, -80.3361269899092, -80.3362524242841, 
    -80.3362747409507, -80.3363932982422, -80.3364158024089, 
    -80.3364967992837, -80.3367162399084, -80.3371325544911, 
    -80.3374427961572, -80.3377270503235, -80.3381239242811, 
    -80.3383631774058, -80.3385746680304, -80.3386230524054, 
    -80.3390010513631, -80.3396368044872, -80.340570175319, 
    -80.3416210524007, -80.3421557357332, -80.3426319836492, 
    -80.3430091773986, -80.3434838596895, -80.3444324930214, -80.34532041802, 
    -80.3453770513532, -80.3458733721858, -80.3464452336433, 
    -80.3471756773921, -80.3478980503077, -80.3481841711405, 
    -80.3488356732229, -80.349427301347, -80.3498942378046, 
    -80.3499584211378, -80.3500224253044, -80.3504314232204, 
    -80.351121111761, -80.3514142325939, -80.3515339878021, 
    -80.3519876096763, -80.3521701763427, -80.3525216784255, 
    -80.3530355482164, -80.3531566107162, -80.353509365924, -80.353903235715, 
    -80.354317608631, -80.3546529909222, -80.3548693617552, 
    -80.3549853596717, -80.3550927971715, -80.355197604463, 
    -80.3552201815463, -80.3552429315463, -80.3553274867544, 
    -80.3554562377959, -80.3559301752952, -80.3563654273779, 
    -80.3569391773769, -80.3573741763346, -80.3581251107084, 
    -80.3584027971664, -80.3585625492494, -80.3588019252907, 
    -80.3590209200821, -80.3591634252902, -80.3593249263316, 
    -80.3594662357063, -80.3596464200811, -80.3597583659143, 
    -80.3600687357055, -80.3603284242467, -80.3605683586213, 
    -80.3608801086208, -80.3613126742452, -80.3615892357031, 
    -80.3620842377857, -80.3627389232013, -80.3628399252845, 
    -80.362927363826, -80.3632118638255, -80.3634706117418, 
    -80.3638474898663, -80.3640867388242, -80.3641164221575, 
    -80.3641222377825, -80.3641393648658, -80.3641517992407, 
    -80.3641790534074, -80.3642421846573, -80.3642908034072, 
    -80.3643054888238, -80.3643981773654, -80.3644649252819, 
    -80.3647733627815, -80.3653731752805, -80.3658529273631, 
    -80.3661956690293, -80.366589802362, -80.3667152367368, -80.367001050278, 
    -80.3674466159023, -80.3677207992353, -80.3679606836099, 
    -80.3681694211095, -80.3685947356922, -80.3691259283997, 
    -80.369571484649, -80.3701712992314, -80.3704282971477, 
    -80.3707024242306, -80.3710772981884, -80.3713413586046, 
    -80.3717537981873, -80.3722266721449, -80.3729344252688, 
    -80.3732874242266, -80.3735016763096, -80.3737359877676, 
    -80.3738089888091, -80.3740306096421, -80.3746818617244, 
    -80.3748995585991, -80.3751171763071, -80.3757504856811, 
    -80.3763633606802, -80.376717800263, -80.3767970502628, 
    -80.3768341106794, -80.3768299273461, -80.3770274221375, 
    -80.3773857950536, -80.3778438638029, -80.3780851773441, 
    -80.3783237388021, -80.3782866763022, -80.378150989844, 
    -80.3781534263024, -80.3782769200522, -80.3783482367188, 
    -80.3784136752603, -80.3787735450514, -80.3792190513007, 
    -80.3796303023418, -80.3800879262994, -80.3802219231741, 
    -80.3807166158817, -80.3814712981722, -80.3815093617138, 
    -80.3820232377547, -80.3823408627542, -80.382515922129, 
    -80.3831324856696, -80.3834190492109, -80.3838107398353, 
    -80.3845902356674, -80.3848904887919, -80.3851054867083, 
    -80.3853712919162, -80.3856604210824, -80.3859488606653, 
    -80.3862584283732, -80.386528674206, -80.3867611752473, 
    -80.3866903669141, -80.3864161762896, -80.3863990492063, 
    -80.3865018627478, -80.3866217992059, -80.3869474210804, 
    -80.3875814221211, -80.3875981137877, -80.3877361117042, 
    -80.3885306752446, -80.388690985661, -80.388699054411, -80.3887328012859, 
    -80.3889711700356, -80.3892359856602, -80.3896891710762, 
    -80.3903917367001, -80.3906830471163, -80.3907858648244, 
    -80.3908591137827, -80.3909059273242, -80.3909743606575, 
    -80.3910429231574, -80.391282863782, -80.3917454887813, 
    -80.3921568012806, -80.392585173155, -80.3930992408625, 
    -80.3933221189872, -80.3934076741954, -80.3935619252368, 
    -80.3936612377366, -80.3939654231528, -80.3944406148187, 
    -80.3944759273187, -80.3948172346098, -80.3957283012751, 
    -80.3965413627321, -80.3976923616887, -80.3986858054372, 
    -80.3993873668944, -80.3994022991861, -80.3996424877274, 
    -80.3997436127272, -80.3998508710604, -80.4000050533518, 
    -80.4001764241848, -80.4003477991846, -80.4005534221009, 
    -80.4007590502256, -80.4009024273087, -80.401365611683, 
    -80.4018990502238, -80.4025720543895, -80.4031067398053, 
    -80.4040361731372, -80.404768738761, -80.4057195523013, 
    -80.4061852387588, -80.4063725502169, -80.4073601752154, 
    -80.407789986673, -80.4080761762559, -80.4083331731305, 
    -80.4085388033386, -80.4087787377132, -80.4091728606292, 
    -80.4097554845866, -80.4100707991695, -80.4101871731277, 
    -80.4105616137521, -80.4109568054181, -80.4112543647927, 
    -80.4112712387509, -80.4115515512505, -80.4118077356251, 
    -80.4120230481248, -80.4123173627077, -80.4127701147903, 
    -80.4134414252059, -80.4149439241619, -80.4157956814523, 
    -80.4164515502013, -80.4173447397832, -80.4180586126988, 
    -80.4186159887396, -80.4189723595724, -80.41937086478, -80.4196129251964, 
    -80.4196514897797, -80.4196963022795, -80.4201158564456, 
    -80.4208697376944, -80.4210482366524, -80.4217203626931, 
    -80.423479738732, -80.4242794866474, -80.4242846793558, 
    -80.4242879262308, -80.4243933647722, -80.4247248043551, 
    -80.4249658637297, -80.4250713637296, -80.4249206783131, 
    -80.4246645491468, -80.4245138626887, -80.4244276803972, 
    -80.4243783012306, -80.4243632366473, -80.4243632418556, 
    -80.4244384876889, -80.4245126137304, -80.4246043022719, 
    -80.4248001741466, -80.4251164866461, -80.4254178647707, 
    -80.4255986772704, -80.425598678312, -80.4255233668538, -80.425432985604, 
    -80.4252822970626, -80.4251918606043, -80.425191871021, -80.425206986646, 
    -80.425237111646, -80.4252521731042, -80.4252672345626, 
    -80.4251316074794, -80.4248754876882, -80.4244536116472, 
    -80.4240124220645, -80.4239413626896, -80.4232633595657, 
    -80.4226305501917, -80.4222238001923, -80.4218320512346, 
    -80.421530676235, -80.4212896126937, -80.4208979272777, 
    -80.4205965512365, -80.4203554856119, -80.4202048626954, 
    -80.4201144293622, -80.4201294845706, -80.4202651064454, 
    -80.4204032397785, -80.4204158001951, -80.4204911116533, 
    -80.4205061710283, -80.4205212293616, -80.4203856095701, 
    -80.4202350543621, -80.4200692376957, -80.4198582991543, 
    -80.4194967387382, -80.4193027262385, -80.4191200491554, 
    -80.4186529845728, -80.4183516783233, -80.4181708637403, 
    -80.4179900491572, -80.4177188606159, -80.4175681710329, 
    -80.417477177283, -80.4174175481164, -80.4173421720749, 
    -80.4171613595752, -80.4169364199922, -80.4168600512423, 
    -80.4164683606179, -80.4164080522847, -80.4164833627012, 
    -80.4166641752009, -80.4171764272835, -80.4174326147831, 
    -80.4177489887409, -80.4180201751988, -80.4183818001983, 
    -80.4184316116565, -80.4187433606144, -80.4190748606139, 
    -80.4191501772804, -80.4191232408221, -80.4191049856138, 
    -80.4189994876973, -80.4188036762393, -80.4185997356146, 
    -80.4185749908229, -80.4180559887404, -80.4171835533251, 
    -80.4168090502007, -80.4167521783258, -80.416611112701, 
    -80.4162948627015, -80.4158510522855, -80.4156518033275, 
    -80.4155088637444, -80.4156602335358, -80.4154279804112, 
    -80.4152862366614, -80.4145397991626, -80.4139371158302, 
    -80.4136208012473, -80.4134851127059, -80.4133061804145, 
    -80.4132289897896, -80.4130481814565, -80.4129879262483, 
    -80.4129879262483, -80.4128824845818, -80.4125961783323, 
    -80.4121442377079, -80.4118579231251, -80.4112703627093, -80.41083342521, 
    -80.4106224866686, -80.4103211741691, -80.409963860628, -80.409929426253, 
    -80.4094322450038, -80.4089049304213, -80.4082721116723, 
    -80.4076242387566, -80.4066448637582, -80.4060121137591, 
    -80.4054997991766, -80.4047766158444, -80.4040835460538, 
    -80.4035110398047, -80.4030741137637, -80.4023961127231, 
    -80.4017030481408, -80.4012661148082, -80.4008141158506, 
    -80.4004014200178, -80.4002286731431, -80.4001993627265, 
    -80.3998046752271, -80.3996991793939, -80.3995636137691, 
    -80.3993376210611, -80.3990814231449, -80.3987499866871, 
    -80.3981774887713, -80.3977984283552, -80.3973939866892, 
    -80.3966561773153, -80.3965050533572, -80.3959624898164, 
    -80.3953836148173, -80.3940130523194, -80.39255923878, -80.3910971148239, 
    -80.3891953658686, -80.3878844242039, -80.3865494200393, 
    -80.3856149887908, -80.3854311085827, -80.3851972387914, 
    -80.3848887377503, -80.3841353648348, -80.3838189887936, 
    -80.3836080481689, -80.3834874908774, -80.3833519252526, 
    -80.383110859628, -80.3828324856701, -80.3827040512953, -80.382236988796, 
    -80.3817849867134, -80.3815138002555, -80.3812878012975, 
    -80.381016613798, -80.3803235471323, -80.3798715429664, 
    -80.3795701710918, -80.3793290481755, -80.3791031148426, 
    -80.3788620471346, -80.3786715471349, -80.3786661710932, 
    -80.378619547135, -80.3784475513019, -80.3783949835936, 
    -80.3781086742191, -80.3777621742196, -80.3774862992201, 
    -80.3773554200536, -80.376873299221, -80.3765267356799, 
    -80.3762404856804, -80.3760596731806, -80.3759089835975, 
    -80.3756227377646, -80.3751104846404, -80.3741661731835, 
    -80.3729201127688, -80.3724097961029, -80.3720261117285, 
    -80.3716488013125, -80.3714685533961, -80.3714569263128, 
    -80.3714463627711, -80.3712240471465, -80.3708632419387, 
    -80.3703063013145, -80.37002736069, -80.3697077388155, -80.3694669242325, 
    -80.369368738816, -80.3693399856911, -80.3688729211084, 
    -80.3685263638173, -80.368315428401, -80.368059291943, -80.36784835861, 
    -80.3676524867353, -80.3674716773606, -80.3671854263194, 
    -80.3667785502784, -80.3664170481956, -80.3662781148625, 
    -80.3658442377798, -80.3655682961136, -80.3652112961141, 
    -80.3646961096566, -80.3645176731985, -80.3639541752827, 
    -80.3638246127829, -80.3637561106997, -80.3635049888251, 
    -80.3631087346591, -80.3627487940346, -80.3623099877853, 
    -80.3621286117439, -80.3619676784108, -80.3618864825776, 
    -80.3615893607031, -80.3611743648704, -80.3606596117462, 
    -80.3601643013303, -80.3598994232057, -80.3598178659142, 
    -80.3593959804982, -80.3593421075816, -80.3591549190402, 
    -80.3587933648741, -80.3585371148745, -80.35816054925, -80.3577838648757, 
    -80.3574373638345, -80.3572414867515, -80.3571510492516, 
    -80.3571050513351, -80.3570733013351, -80.3569913627936, 
    -80.3567717982106, -80.3564942377943, -80.3559802971701, 
    -80.3553887357127, -80.3547590523804, -80.354093175298, 
    -80.3542530534228, -80.3543140492561, -80.3543134909227, 
    -80.3542968013394, -80.3542988002977, -80.3542413627978, 
    -80.3540451127981, -80.3538102930068, -80.3535747919655, 
    -80.3532796127993, -80.3530818575913, -80.3527836128001, 
    -80.3525659253004, -80.352151612801, -80.3518948607181, 
    -80.3516178607185, -80.3512131805109, -80.3510815482194, 
    -80.3505462398869, -80.3497150513465, -80.3492795503055, 
    -80.3489029888478, -80.3486871680147, -80.3485315471817, 
    -80.3484479888485, -80.3481782982239, -80.3479811763492, 
    -80.3476649273913, -80.3474272992667, -80.3471687398921, 
    -80.3465760534347, -80.3461051128104, -80.3456980503111, 
    -80.3455373659363, -80.3451396107286, -80.3443081784382, 
    -80.343812797189, -80.3437812992724, -80.3432956836481, 
    -80.3430559836485, -80.3429536128153, -80.3428329242739, 
    -80.3424784867744, -80.3413337982345, -80.3411836096931, 
    -80.3409858003184, -80.3405084274025, -80.3404688013609, 
    -80.3402090482363, -80.33991173782, -80.3391594878212, -80.3390292409464, 
    -80.3390259253214, -80.3388451784467, -80.3387095513636, 
    -80.338483545114, -80.3383866732391, -80.3382876794893, 
    -80.3381458607395, -80.3380767399062, -80.3378356711566, 
    -80.3376548607403, -80.3374741086572, -80.3373084211574, 
    -80.337172738866, -80.3369166096997, -80.3367876701166, 
    -80.3361479284509, -80.3357517399099, -80.3357323586599, 
    -80.3357125513683, -80.3357890472014, -80.33562998991, -80.3351949263691, 
    -80.3344022326203, -80.3340901784541, -80.3339073649127, 
    -80.3333129263719, -80.3323994867901, -80.331824296166, 
    -80.3316739867912, -80.3315247388747, -80.3309972378339, 
    -80.330710613876, -80.3301546117935, -80.3296196086694, 
    -80.3294208617947, -80.3292032378367, -80.3287101107541, 
    -80.3285007420045, -80.3284925482545, -80.3284749232545, 
    -80.3282345513799, -80.3281936701299, -80.328127735755, 
    -80.3279316815887, -80.3277709232556, -80.3272736753397, 
    -80.327251364923, -80.3266697982573, -80.3264302367993, 
    -80.3261590503414, -80.3261289867998, -80.3260837357582, 
    -80.3260686763832, -80.3260936784665, -80.3260987972165, 
    -80.326174113883, -80.3262946763829, -80.3263097367995, 
    -80.3261289222165, -80.3257221086754, -80.3251496138847, 
    -80.3248181118018, -80.3246373586771, -80.324516800344, 
    -80.3244264253441, -80.3241877378445, -80.3237189847202, 
    -80.3231868576377, -80.3224754868055, -80.3219584222229, 
    -80.3219224263897, -80.3214482399321, -80.3209939857661, 
    -80.3204346743086, -80.3199992357676, -80.3194423013935, 
    -80.3193116743104, -80.3190749878524, -80.3188381784778, 
    -80.3184523003534, -80.3182851722286, -80.3180493618123, 
    -80.3179932441041, -80.3179716784791, -80.3178990493126, 
    -80.3178426753543, -80.3177859243127, -80.3175891170214, 
    -80.3172533586886, -80.3168244878559, -80.316799053481, 
    -80.3167862388976, -80.3166406107729, -80.3166023638979, 
    -80.3165257993147, -80.3164569899398, -80.3164088628565, 
    -80.316363174315, -80.3161132368153, -80.316094984732, -80.3158186107741, 
    -80.3156516774411, -80.3151371139002, -80.3147226805675, 
    -80.3143084253598, -80.3134604222361, -80.3131289826533, 
    -80.312657298279, -80.3121344889049, -80.31202579828, -80.3114618618226, 
    -80.3111158024481, -80.3107002316154, -80.3106858691154, 
    -80.3106189232822, -80.3104204889075, -80.3101044909913, 
    -80.3099261066166, -80.3098286701584, -80.309671675367, 
    -80.3094154889091, -80.309269736826, -80.3092633628676, 
    -80.3091002993262, -80.3087871774517, -80.3084542316189, 
    -80.3080426128695, -80.3075678618286, -80.3066862347466, 
    -80.3063697993305, -80.3061417368308, -80.3057973607897, 
    -80.3049359878743, -80.3043332378753, -80.3041049847507, 
    -80.3039949180841, -80.3037814868345, -80.3034474253767, 
    -80.3028523639193, -80.302564047253, -80.3021640545453, 
    -80.3017816128793, -80.3013501087133, -80.300888927464, 
    -80.3003831701731, -80.2996481722575, -80.2994696753829, 
    -80.2993930482996, -80.2994352982996, -80.2992791076748, 
    -80.2991619847583, -80.2991833014249, -80.2991061128834, 
    -80.2989109878837, -80.2985371160093, -80.2982070483015, 
    -80.2973718618445, -80.2969657368451, -80.2968399222619, 
    -80.2967544253871, -80.2965039889291, -80.2960482983048, 
    -80.2957914243469, -80.2957557972636, -80.2956559910137, 
    -80.2956547045554, -80.2956169858055, -80.2957700524719, 
    -80.2957036170553, -80.2956602347638, -80.2955676108056, 
    -80.2952737972644, -80.2951572399729, -80.2949627368482, -80.29487417539, 
    -80.2948423618483, -80.2946088628904, -80.2943006097659, 
    -80.2940026160163, -80.2937436139334, -80.2933659941423, 
    -80.2924216753938, -80.2920170493528, -80.2916232993534, 
    -80.2914754201869, -80.2912933024789, -80.2912516753956, 
    -80.2910471774792, -80.2908646128962, -80.2907516743547, 
    -80.2907390535214, -80.2907096108131, -80.2907137941464, 
    -80.2907845503963, -80.2910933639375, -80.2913296774788, 
    -80.2913681743537, -80.291458982687, -80.2917096139366, 
    -80.2917977972697, -80.2915783576868, -80.2916899837282, 
    -80.2917980524781, -80.2920735472693, -80.2925067389353, 
    -80.2930003024762, -80.2933219847674, -80.2933948056006, 
    -80.2936501139336, -80.2941236733078, -80.2941624233077, 
    -80.2940221160163, -80.2938616722665, -80.2939372378914, 
    -80.2940726108079, -80.2941499941411, -80.2941897993493, 
    -80.2944884253906, -80.2945661764321, -80.2944835514322, 
    -80.2944552410156, -80.2945059868489, -80.2944847378906, 
    -80.2943646753907, -80.2940865524745, -80.2943794889324, 
    -80.294673798307, -80.2951067347646, -80.2955778014306, 
    -80.2958505483051, -80.2959107399717, -80.2959862368466, 
    -80.295908860805, -80.2958605493468, -80.2958988003884, -80.296135300388, 
    -80.2964373024709, -80.2965108618458, -80.2968339264286, -80.2970522951783 ;

 y = 36.5354153651647, 36.5357538641225, 36.5360843026637, 36.5363068641217, 
    36.5364974912047, 36.536740801621, 36.5367946745376, 36.5371058016204, 
    36.5374752422449, 36.5379336151608, 36.5382661828686, 36.5386683037013, 
    36.5389823026592, 36.5391110547423, 36.5390962391173, 36.5390719912007, 
    36.5388839266176, 36.5383971141184, 36.5379323057858, 36.5375498037031, 
    36.5373198641201, 36.5369536172457, 36.5363746755799, 36.5361129912053, 
    36.5358550537057, 36.5356335557894, 36.5354722412063, 36.5353808037064, 
    36.5353074922482, 36.5353897391231, 36.5356388641227, 36.5357619266225, 
    36.5358607380807, 36.5360088630804, 36.5359395505806, 36.5358165505808, 
    36.5355549870395, 36.5353544287065, 36.5351259307902, 36.5349533026654, 
    36.5349404870404, 36.5348146193323, 36.5346784287075, 36.5344878037078, 
    36.5344187401662, 36.5345089912078, 36.5346238641243, 36.5346417995409, 
    36.5346480526659, 36.5346543016242, 36.5348969912072, 36.5351281807901, 
    36.5352634891233, 36.5353703641231, 36.5355057422479, 36.5355530537062, 
    36.5357417432892, 36.5358834912057, 36.5360676182887, 36.5361331172469, 
    36.5360221141221, 36.5359723037055, 36.5356732432893, 36.5354138005814, 
    36.53523268079, 36.5351029953735, 36.535031931832, 36.5348527995406, 
    36.534590177666, 36.5342861162081, 36.5340398037085, 36.5338600568338, 
    36.533695800584, 36.5336773630841, 36.5335453026676, 36.5333843703762, 
    36.5332259880848, 36.5330869297517, 36.5328199912104, 36.5327476787105, 
    36.5326211141274, 36.5325685505858, 36.5325171172526, 36.532429619336, 
    36.5321458026698, 36.53200411517, 36.5320691755866, 36.5321057412115, 
    36.5323289922528, 36.5324073026694, 36.5324285526693, 36.5324301172527, 
    36.5325178662109, 36.5326246755857, 36.5328457401687, 36.5331133672516, 
    36.5331527412099, 36.5334522412094, 36.533718616209, 36.5338444901672, 
    36.5339744307919, 36.5340340495419, 36.53417511725, 36.534604049541, 
    36.5346849255825, 36.5346989287075, 36.5346531172492, 36.5345494922494, 
    36.5343978016246, 36.5342559891249, 36.5342000526666, 36.5342110516249, 
    36.5342214901665, 36.5342128005833, 36.5340986776667, 36.533917427667, 
    36.5337266797507, 36.533724363084, 36.5334790526677, 36.5333239255846, 
    36.5332394266264, 36.5330539297517, 36.5330291766268, 36.5328176162104, 
    36.5323747422528, 36.5320656120449, 36.5319144901702, 36.5317719235037, 
    36.5314209266293, 36.5311823662129, 36.5309154901717, 36.5306406162138, 
    36.5303464276726, 36.5300425505897, 36.5296734912153, 36.5294638005906, 
    36.5294698672573, 36.5294740526739, 36.5295613057988, 36.5295719880904, 
    36.5295062422572, 36.5293454297575, 36.5292471172576, 36.5291468026745, 
    36.5289671745497, 36.5287248016334, 36.5286561141335, 36.5284353037172, 
    36.5284150547589, 36.5281423037177, 36.5281916172593, 36.5282529901758, 
    36.5284118026756, 36.5286800537168, 36.5289006818415, 36.5291212380911, 
    36.5292941172576, 36.5295436703822, 36.5298120516317, 36.5302004912145, 
    36.5307969964219, 36.5311499932963, 36.5314453610042, 36.5316646162122, 
    36.5319224287118, 36.5322120537114, 36.5323539287111, 36.5325372391275, 
    36.532635121419, 36.532675302669, 36.5327341172522, 36.5328395526687, 
    36.5329922370435, 36.5333548047512, 36.5336699880841, 36.5337461182923, 
    36.5340991776667, 36.5343188651664, 36.5345198651661, 36.5347601141241, 
    36.5349913057904, 36.5351262995401, 36.5352038037067, 36.5353864964147, 
    36.5355398047478, 36.5356741141226, 36.5357419255809, 36.5358308651641, 
    36.5359669276639, 36.5361603672469, 36.5364388641215, 36.5365530537046, 
    36.536522299538, 36.5363636141216, 36.5361093026636, 36.5358067380808, 
    36.5355995526644, 36.5354556182896, 36.535247427665, 36.5350554932903, 
    36.5348799287072, 36.5347251120408, 36.5347050547492, 36.5345933016243, 
    36.5346577401659, 36.5348126818323, 36.5350059870403, 36.5350929287069, 
    36.5351608026651, 36.5351138005818, 36.5349234912071, 36.5346853651658, 
    36.5346293099576, 36.5344575516245, 36.5342297391249, 36.5338404891255, 
    36.5334792401677, 36.5333749922512, 36.5332905485013, 36.5332453651681, 
    36.5331859912098, 36.5331810547515, 36.533078056835, 36.532850929752, 
    36.5326042391274, 36.5320918682949, 36.5318835474619, 36.5317328016288, 
    36.5316501787122, 36.5316909349622, 36.5317407401704, 36.5317034912121, 
    36.5316084891289, 36.5314172401709, 36.5310254901715, 36.5305194245473, 
    36.5302385526728, 36.530043740173, 36.5298350516317, 36.5294555547573, 
    36.5292850516325, 36.5292571120493, 36.5292886172576, 36.5293478641324, 
    36.5293977380907, 36.529418802674, 36.5293624932991, 36.5292298016327, 
    36.5290679266329, 36.5288011755916, 36.5285345526754, 36.5282684912175, 
    36.5279930537179, 36.5278135547599, 36.5277298620516, 36.5277751787182, 
    36.5266074901784, 36.5257634901797, 36.5253085516387, 36.5246324287231, 
    36.5239328641409, 36.5237589266411, 36.523637302683, 36.5235469870581, 
    36.5233429266418, 36.5231679891421, 36.522795113101, 36.5222938047684, 
    36.5222412391435, 36.5216588631027, 36.5209119266456, 36.5204450568546, 
    36.520406118313, 36.5200603651886, 36.5194582422728, 36.5190644287318, 
    36.5186234276908, 36.5181939912331, 36.5178436141503, 36.5175804933174, 
    36.5167732412353, 36.5157707412369, 36.5152942412376, 36.5149058058216, 
    36.5147034901968, 36.5146799881136, 36.5144454287389, 36.5142639266559, 
    36.514197492281, 36.5140339276979, 36.5136855516567, 36.5134911766571, 
    36.5131578672826, 36.5129764901995, 36.5127103631166, 36.5125938662418, 
    36.5124903027003, 36.5121592422842, 36.5117310537431, 36.5110684245775, 
    36.5106250506199, 36.5107927995779, 36.5111869266606, 36.5112896162438, 
    36.5112056777023, 36.5111631183274, 36.5110700527025, 36.5109947391609, 
    36.5109344912444, 36.5108139256196, 36.5106934277031, 36.5104221787452, 
    36.510344926662, 36.5100304922875, 36.5097140527046, 36.5094127422884, 
    36.509253306872, 36.509021301664, 36.5083579297901, 36.5082751224985, 
    36.5081406787487, 36.5078929256241, 36.5073651766666, 36.507130489167, 
    36.5069973662505, 36.5067300485426, 36.5067262412509, 36.5067271787509, 
    36.5066265547927, 36.5064233027097, 36.506256180835, 36.5060464891686, 
    36.5057016131275, 36.5054459891696, 36.5051689902116, 36.5049121141704, 
    36.5047470547956, 36.5047046141707, 36.5048663662538, 36.5049874902119, 
    36.5046856766708, 36.5047068620873, 36.5043688037546, 36.5042901162547, 
    36.5043467422963, 36.504336677713, 36.5043804881295, 36.5043202422963, 
    36.5041846152132, 36.5040188683384, 36.5039668631302, 36.5039284922969, 
    36.5039586110469, 36.5040490527134, 36.5042298037548, 36.5043804891712, 
    36.5044859912544, 36.5045010527127, 36.5044256777128, 36.5042298068798, 
    36.5040339297968, 36.5038629277137, 36.5038230537554, 36.5035518006308, 
    36.5032956797979, 36.5032446787563, 36.5031299891731, 36.5030071162567, 
    36.5029492422984, 36.5029492402151, 36.502994365215, 36.5029943662567, 
    36.5029039912569, 36.5027382422988, 36.5025122412574, 36.5021204881331, 
    36.5018493016751, 36.5015781152172, 36.5012767975094, 36.5010055589681, 
    36.500659054802, 36.5003577423025, 36.5001640527194, 36.4999057412615, 
    36.4996834902201, 36.4993331777207, 36.4991401162627, 36.498472740222, 
    36.4982123027224, 36.4980024902228, 36.4981493641809, 36.498307810014, 
    36.4984131798055, 36.4985457370969, 36.4985705506386, 36.4985949287635, 
    36.4986099902218, 36.4986551787634, 36.4987606766799, 36.4989414277213, 
    36.4990079245962, 36.4989405527213, 36.4988818662631, 36.4990774245961, 
    36.499132555846, 36.4993003652208, 36.4994044902206, 36.4994537412622, 
    36.4994537412622, 36.499378367304, 36.4991523631377, 36.4988811787631, 
    36.4986400516801, 36.498504549597, 36.4984743641804, 36.4984743620971, 
    36.4984894287637, 36.4987455537633, 36.4988265548049, 36.4989715485546, 
    36.4990921120961, 36.4991222370961, 36.4990600527211, 36.4989866829296, 
    36.4988811808464, 36.4988617402215, 36.4988510527215, 36.4988811766797, 
    36.4987757412633, 36.4986702412634, 36.4983688652222, 36.4981929923058, 
    36.4980073037644, 36.497675866265, 36.4974950516819, 36.4972991798072, 
    36.4970882412659, 36.4969526745994, 36.4967718693914, 36.4967534214747, 
    36.4965157423084, 36.4963499891837, 36.4962143662672, 36.496093864184, 
    36.4959130516843, 36.4955966777265, 36.4955368662683, 36.4955092381433, 
    36.495473301685, 36.495281365227, 36.4950727402273, 36.4947177402279, 
    36.4945391777281, 36.4942336798119, 36.4938810516875, 36.493575614188, 
    36.4934069277299, 36.4933065496051, 36.4930654923138, 36.4927339881476, 
    36.4923724246065, 36.4919053641906, 36.4912876141915, 36.4908657381505, 
    36.4905794860676, 36.4902329266932, 36.4898412402354, 36.4894494256527, 
    36.4891782350281, 36.4889372371118, 36.4885605548208, 36.4883836121127, 
    36.4881386766965, 36.4878072412803, 36.4875360496141, 36.487129242323, 
    36.4869183048233, 36.4865717371155, 36.4863306777409, 36.486029366283, 
    36.4858033642, 36.4856526787836, 36.4855773642004, 36.4854417433673, 
    36.485438491284, 36.4852006777426, 36.4848843037848, 36.4845829871186, 
    36.4842665496191, 36.483920054828, 36.483694052745, 36.4833625558705, 
    36.4829859256628, 36.4824585548303, 36.4821890527473, 36.4819764277477, 
    36.4816148006649, 36.4813587392069, 36.4811628673323, 36.4809519298326, 
    36.4806204298331, 36.4803341767085, 36.4801081777505, 36.4799273631675, 
    36.4797616756678, 36.4794000527517, 36.4790384277522, 36.4786015517112, 
    36.4783906142115, 36.4782248662951, 36.4780289892121, 36.4778933662956, 
    36.4778029871291, 36.4776891777543, 36.4775920537961, 36.477456492338, 
    36.4772606162966, 36.4767935506724, 36.4764319277563, 36.4761004902568, 
    36.4754375537995, 36.474880051717, 36.4744733017176, 36.4741267381765, 
    36.4740659298433, 36.4739158642185, 36.4737500496354, 36.4735240517191, 
    36.4732829902612, 36.4730720548448, 36.4728913017201, 36.4727899256786, 
    36.4725447392206, 36.4720475517214, 36.4714147381807, 36.4713056152642, 
    36.4711702381811, 36.4697061111, 36.4689994892261, 36.4682815496439, 
    36.4682483642273, 36.4680247402693, 36.4677686152697, 36.4673919902703, 
    36.4671358027707, 36.4668495517295, 36.4665783673549, 36.4663222402719, 
    36.4660752423557, 36.4660058642308, 36.4656593038147, 36.4653579881901, 
    36.4647552975661, 36.4641224934004, 36.4636704913177, 36.4631883652768, 
    36.4630703038187, 36.4627664881941, 36.462450115278, 36.4621036173618, 
    36.4617419975708, 36.4614822423628, 36.4610489225718, 36.4606421111141, 
    36.4602051809064, 36.4599189298652, 36.4595874913241, 36.4593011798662, 
    36.4591053027831, 36.4589244882001, 36.4586684267422, 36.4585328048674, 
    36.4583068007011, 36.4579301132017, 36.4575986736188, 36.4571768017445, 
    36.4568989288283, 36.4567247986202, 36.4561221163294, 36.4557906809133, 
    36.4554441184138, 36.4551729267476, 36.4550223038312, 36.4547812382065, 
    36.4545939892485, 36.4544648017487, 36.4541785569575, 36.4539676142495, 
    36.4538466152913, 36.4537265507082, 36.4536210527917, 36.4535758632084, 
    36.4535156173752, 36.4533197402922, 36.4531691152924, 36.4530184277926, 
    36.452973236126, 36.4528526152928, 36.4526718652932, 36.4524609267518, 
    36.4522198663355, 36.4518281767528, 36.4513158652953, 36.4510296184207, 
    36.4509221194625, 36.4506228017547, 36.4502913663385, 36.4500205538389, 
    36.450003803839, 36.4498876767558, 36.4498294298809, 36.4495289892564, 
    36.449137239257, 36.448670178841, 36.4483688048832, 36.4480524892587, 
    36.4476155517593, 36.4470731194685, 36.4468621767605, 36.446560867386, 
    36.4462321757198, 36.4461389903033, 36.4456869913457, 36.4453555538462, 
    36.4451069319716, 36.4448056173887, 36.4445645517641, 36.4443084267645, 
    36.4439618653067, 36.4436003028072, 36.4432537434328, 36.443103052808, 
    36.4430729246831, 36.4431784288495, 36.4433441778076, 36.4435744330156, 
    36.4436153642656, 36.4438865507234, 36.4441124882231, 36.4442330528062, 
    36.4442782986395, 36.4442933653061, 36.444202928848, 36.4440070528066, 
    36.4438413038485, 36.4436153642656, 36.4435249278073, 36.4433893642659, 
    36.4431633028079, 36.4428017403085, 36.4427749278085, 36.4425305507256, 
    36.4424099913508, 36.4423982434341, 36.4423648028092, 36.4423798642674, 
    36.4424099923924, 36.4423949278091, 36.4423045517676, 36.4419579903098, 
    36.4416416142686, 36.4415362444771, 36.4412951121858, 36.4411370496861, 
    36.4411336788527, 36.4410546767695, 36.4409982330196, 36.4410454892695, 
    36.4410580517695, 36.4414058653106, 36.4419789278097, 36.4422875517676, 
    36.4425536788505, 36.4431914882245, 36.4436049319739, 36.4438212413485, 
    36.4441596142647, 36.4444437403059, 36.4448866757219, 36.4453308028046, 
    36.4455343028042, 36.4454949871793, 36.4453638038461, 36.4450900528049, 
    36.4447851163471, 36.4444964288475, 36.444383365306, 36.4444573028059, 
    36.4444617434309, 36.444588114264, 36.4445541767641, 36.4443926163477, 
    36.4442755548895, 36.4441138007231, 36.4438224944735, 36.4433941173909, 
    36.4430513632248, 36.4427258028086, 36.4423316778092, 36.4420168590597, 
    36.4417106778101, 36.4415779267687, 36.4415953048937, 36.4416386173936, 
    36.4418734934349, 36.4419976163514, 36.4420089913514, 36.4421181142679, 
    36.4422106153094, 36.4421599923928, 36.4419834288514, 36.4418861215599, 
    36.4415776778104, 36.4411835548943, 36.4411664298943, 36.4413549288524, 
    36.4418176142683, 36.4423076798926, 36.4425347382256, 36.4429169903083, 
    36.4429295517666, 36.4435204278074, 36.4441384944731, 36.4446758017639, 
    36.4449753017634, 36.4451623673881, 36.4452765538463, 36.4452882392629, 
    36.4453657403045, 36.4453051153046, 36.4452619913463, 36.4450391757217, 
    36.4447135538472, 36.4446793017639, 36.4446793059305, 36.4448335528053, 
    36.4449706194717, 36.4450734278049, 36.4451419882215, 36.445296176763, 
    36.4457417434289, 36.4459286153036, 36.4462215590531, 36.4464100528029, 
    36.446547117386, 36.4466499267608, 36.4467017340524, 36.4468100507189, 
    36.446952612177, 36.4471846132183, 36.4472399267599, 36.4475106153012, 
    36.4479699309255, 36.4480473028003, 36.4480551153003, 36.4483293080082, 
    36.4485863048828, 36.4489290548823, 36.4494259871732, 36.4498029892559, 
    36.4502313642553, 36.4504319923799, 36.4506316767547, 36.4507266788378, 
    36.450835552796, 36.4508676777959, 36.4508602361293, 36.4508256767543, 
    36.4507759892544, 36.4507209288378, 36.4506678642546, 36.450627675713, 
    36.4505723663381, 36.4504352444633, 36.4503605517551, 36.4502249892553, 
    36.4501903642553, 36.4502009288386, 36.4504099288383, 36.4504553027966, 
    36.4504972382132, 36.4505055538382, 36.4505398017548, 36.4507797402961, 
    36.4511053007122, 36.4512897402953, 36.4513398038369, 36.4519463017526, 
    36.4522498017521, 36.4527648038347, 36.4529056777928, 36.4530641757092, 
    36.4535581809168, 36.4539711757078, 36.4542728038323, 36.454239864249, 
    36.4537126163332, 36.4536208027916, 36.4534244892503, 36.4532309277923, 
    36.4532117402923, 36.4532723652922, 36.4532871777922, 36.4533019934171, 
    36.4531388642508, 36.4529574257094, 36.4528976777928, 36.4525130527934, 
    36.4521124923774, 36.4517432423779, 36.451228300712, 36.4510021142541, 
    36.4506644892546, 36.4504753652965, 36.4500599902972, 36.4497344298811, 
    36.4496144902979, 36.4494773663397, 36.4494088652982, 36.4494946163397, 
    36.4495174913397, 36.449528802798, 36.4495288048814, 36.4494431194648, 
    36.4492203652985, 36.4490416777988, 36.4489633059239, 36.4487748017575, 
    36.4486377465494, 36.448671991341, 36.448894743424, 36.4490831777987, 
    36.4492046798819, 36.4492648673818, 36.4492744267567, 36.4493060548817, 
    36.4495270538397, 36.4496223038395, 36.4496658652978, 36.4501456777971, 
    36.4501842392553, 36.4503224892551, 36.4505608632131, 36.4507026173795, 
    36.4509089246709, 36.4518499882111, 36.4528719288345, 36.4531270548758, 
    36.4533791194587, 36.4534563673753, 36.4534229330003, 36.4534121142503, 
    36.4534779288335, 36.4535584902918, 36.4536866777916, 36.4539442402912, 
    36.4540370538327, 36.4543076777906, 36.454658362165, 36.4550569267478, 
    36.4555513694553, 36.4557259257051, 36.4559802382047, 36.456171114246, 
    36.4562654871626, 36.456197554871, 36.4561951819543, 36.4562240527876, 
    36.4562376777876, 36.4561553059127, 36.4560933027878, 36.456027802788, 
    36.4560101767463, 36.455980927788, 36.4558448652882, 36.4557053673718, 
    36.4553852423722, 36.4552403027892, 36.4551426142476, 36.4550445548728, 
    36.4548346777898, 36.4547614298733, 36.4547363007066, 36.4547015548733, 
    36.4547101788316, 36.454714680915, 36.4545683684152, 36.4544842996654, 
    36.4542785538323, 36.4539872392494, 36.4538193048747, 36.4537929902914, 
    36.4537521163331, 36.4534546142502, 36.4532596757089, 36.4531283017508, 
    36.4531267382091, 36.4531228048758, 36.4529749902927, 36.4527801788346, 
    36.4526914330015, 36.4526813017515, 36.4524527382101, 36.4523836767519, 
    36.4523969892519, 36.4525706777933, 36.452759743418, 36.4528526163346, 
    36.453182366334, 36.4536404871666, 36.4539883642494, 36.4542579288324, 
    36.4543200517489, 36.4545919361235, 36.4548143038315, 36.4549718652896, 
    36.4550389882061, 36.455112363206, 36.4552378048725, 36.4554602402888, 
    36.4556834892468, 36.4560028642463, 36.4562441746626, 36.4562896184125, 
    36.4564049309124, 36.4565278017455, 36.45686149237, 36.4570032402864, 
    36.4571111767446, 36.4571306767446, 36.4571391725779, 36.4571034298696, 
    36.4569581152865, 36.4567655517451, 36.456617490287, 36.4564929298705, 
    36.4562008069543, 36.4555044871638, 36.4554904913304, 36.455135616331, 
    36.454891426748, 36.4548455517481, 36.45469724029, 36.4544870527903, 
    36.4544372434154, 36.4545315507069, 36.4546010538318, 36.4546010517485, 
    36.4545668038319, 36.454481116332, 36.4544982434153, 36.454477178832, 
    36.4545164267486, 36.4544824892487, 36.4544836777903, 36.4545124902903, 
    36.4546702413317, 36.4549267413313, 36.4553550548723, 36.4557321152884, 
    36.4560062392463, 36.4560949882045, 36.4561947402877, 36.4563832382041, 
    36.4566231111203, 36.4570343048697, 36.4573771142442, 36.4575869892439, 
    36.4575998673688, 36.4576098642438, 36.4576855548687, 36.4576513048688, 
    36.4576381788271, 36.4575754277855, 36.4573990538275, 36.4571321132029, 
    36.4570933027863, 36.4569311767449, 36.4568026757034, 36.4566418048703, 
    36.4565419267454, 36.4565256788288, 36.4567430527868, 36.4569486798698, 
    36.457239990286, 36.4573942413275, 36.4573429267442, 36.457051553828, 
    36.4566916777869, 36.4564378621623, 36.4564003017457, 36.4559032996631, 
    36.4555987444553, 36.4553703017473, 36.4553702444556, 36.4553039288307, 
    36.4553169277891, 36.4554096132056, 36.4553274913307, 36.4552146132058, 
    36.4550478632061, 36.454902486123, 36.454517797582, 36.4543093673739, 
    36.4538813632079, 36.4536071777917, 36.4533159277921, 36.4530074246676, 
    36.4527846809179, 36.4524590527935, 36.4519449902943, 36.451670801753, 
    36.4514137361284, 36.4513281184202, 36.4513109277952, 36.4512833642536, 
    36.4512260559204, 36.4512558027953, 36.451244175712, 36.4511166798789, 
    36.4507498017545, 36.4502381767552, 36.4498592434225, 36.44931367884, 
    36.4488510517574, 36.4481968028001, 36.4473851142597, 36.4468328642606, 
    36.4465970538442, 36.4466088642609, 36.4466793038441, 36.4468555475938, 
    36.4470440528019, 36.4470440507185, 36.4468384257189, 36.4468069903023, 
    36.4466156798859, 36.446547117386, 36.4465641757193, 36.4465814278026, 
    36.4467527392607, 36.4469926757186, 36.44718117676, 36.447403928843, 
    36.4476950528008, 36.4477123663425, 36.4479865528004, 36.4482023642584, 
    36.4486303611328, 36.448883737174, 36.4486769277993, 36.4483820538414, 
    36.4480187434253, 36.4476439288426, 36.4473000569682, 36.4471104278018, 
    36.4470129278019, 36.4473351153014, 36.4475548632178, 36.447812867384, 
    36.4480659892586, 36.4480753642586, 36.4482240548834, 36.4482592403, 
    36.4481516173835, 36.4479370538422, 36.4477038017592, 36.4476814236342, 
    36.4479226194672, 36.4481553069668, 36.4481546757168, 36.4481543048835, 
    36.4481542361335, 36.4479900496754, 36.4477161142592, 36.4472323048849, 
    36.4469001132188, 36.4463193632197, 36.446108116345, 36.4460354267618, 
    36.4460421673868, 36.4461515538449, 36.4463799298862, 36.4463762100946, 
    36.4463813944696, 36.4466800100941, 36.446779741344, 36.4470826788435, 
    36.4476536757176, 36.4486748027994, 36.4489591142573, 36.4495028632147, 
    36.4501089944638, 36.4504929913382, 36.451021926754, 36.4517437413363, 
    36.452321489252, 36.4527877402929, 36.4531086152925, 36.453381177792, 
    36.4537673673748, 36.454041427791, 36.454250114249, 36.4545863663319, 
    36.454907364248, 36.455357674664, 36.4556795517468, 36.4559678632047, 
    36.4561437434127, 36.4565433027871, 36.4567676767451, 36.4568648027866, 
    36.4569317402865, 36.4569498694532, 36.4570146767447, 36.4572241163277, 
    36.4573714257025, 36.4576131163271, 36.4579493059099, 36.4582060548679, 
    36.4582211163262, 36.4584143017426, 36.4586686163255, 36.4588759309085, 
    36.4591162392415, 36.459197802783, 36.4592449277829, 36.4592449277829, 
    36.4592449298663, 36.459416304866, 36.4597418673655, 36.4602993663229, 
    36.4605473048642, 36.4609756788219, 36.4611214850717, 36.4615754309043, 
    36.4621580506951, 36.4626207392361, 36.4629806809021, 36.4633061777766, 
    36.4638031173592, 36.4641286777754, 36.4644714288165, 36.4647627423577, 
    36.4649169881908, 36.465036927774, 36.4653968631901, 36.4656709308979, 
    36.4657566142312, 36.465834426731, 36.4658594288143, 36.4659794236058, 
    36.4662021798555, 36.4664078048552, 36.4666476756881, 36.4668361788128, 
    36.4670641131875, 36.4672696788122, 36.4675268038117, 36.4677495496447, 
    36.4679551767277, 36.4683664319355, 36.46864061631, 36.468863365268, 
    36.4689319267262, 36.4689661788095, 36.4689661788095, 36.4689545548512, 
    36.4689490517262, 36.4689148017263, 36.4689148017263, 36.4689661788095, 
    36.4691032975593, 36.4691788631842, 36.4693431808923, 36.469497427767, 
    36.4696516808918, 36.4698229881832, 36.4701314892244, 36.4702590538075, 
    36.4720985506797, 36.4724017392209, 36.4726676142204, 36.4730617413032, 
    36.4734729944275, 36.4738499881769, 36.4740041798433, 36.4741584277598, 
    36.4744839913009, 36.4748438642171, 36.4752037381749, 36.4754607402577, 
    36.475769241299, 36.4759405537987, 36.4761119308818, 36.4763346787981, 
    36.4765060517145, 36.4765664267144, 36.4767459881725, 36.4767973652557, 
    36.4769516142138, 36.4772771808799, 36.4776199298378, 36.4779626142122, 
    36.4781168652536, 36.4783738673366, 36.4784912412947, 36.4785966808779, 
    36.4787679902527, 36.4790250475439, 36.4793334923351, 36.4795219923348, 
    36.4797104902512, 36.4797471131678, 36.4799504267091, 36.4799951767091, 
    36.4801731746255, 36.4804130517084, 36.4805330506666, 36.4806358652497, 
    36.4807448037913, 36.4808243631661, 36.4809443027493, 36.4810985517074, 
    36.4813384256653, 36.4815440517066, 36.4818182412895, 36.4819151173311, 
    36.4821438069141, 36.4826064902467, 36.4828806787879, 36.483069183996, 
    36.4831205506625, 36.483034868371, 36.4829663642045, 36.4828978037879, 
    36.4828121110797, 36.4827264298298, 36.4825551142051, 36.4824256142053, 
    36.4822368017056, 36.4820196798309, 36.4820326162892, 36.4822316787889, 
    36.4822455517055, 36.4825839277467, 36.4828709933713, 36.4831731756624, 
    36.4834903652453, 36.4837295548282, 36.4840975579527, 36.4841447423276, 
    36.4842446787858, 36.4846902423268, 36.4849986798263, 36.4853414267008, 
    36.4855299267005, 36.4856841183669, 36.4859411798248, 36.4862324860744, 
    36.4866094871155, 36.4867065516987, 36.4868664912817, 36.4869693006566, 
    36.4871235475313, 36.4873291766977, 36.4873877412809, 36.4874491173225, 
    36.4875176819057, 36.4876204902389, 36.48798036628, 36.4883230516961, 
    36.4886315527373, 36.4889571131535, 36.4892141756531, 36.4894539891944, 
    36.4895775527359, 36.4899408641936, 36.4902131131515, 36.4904999923178, 
    36.4908193037756, 36.4909393641921, 36.4910980506502, 36.4912432402332, 
    36.4915307412745, 36.4917058673159, 36.4918004912741, 36.491821491274, 
    36.491829616274, 36.4919538714822, 36.4922233641901, 36.4925897391895, 
    36.4929726787723, 36.4932924891884, 36.4935954277296, 36.4938818652292, 
    36.494232614187, 36.4944724912699, 36.4947291787695, 36.4949854933525, 
    36.4952409277271, 36.4954809308517, 36.4959943641842, 36.4964763006418, 
    36.496975113141, 36.4972147412657, 36.4975694912651, 36.4978263027231, 
    36.4980985527226, 36.4981409245976, 36.4983544933472, 36.4986629266801, 
    36.498937116263, 36.499125615221, 36.4992113027209, 36.4993484287623, 
    36.499605428762, 36.4997939287617, 36.4998967391782, 36.4998967412615, 
    36.4998281787616, 36.4997768016784, 36.4997253662618, 36.4996397391786, 
    36.4993792391789, 36.499348426679, 36.4990056777212, 36.4989199902213, 
    36.4990056777212, 36.4992112985543, 36.4994512433455, 36.4996137423036, 
    36.4996293620953, 36.499536181887, 36.4993783037623, 36.499367176679, 
    36.4997082412618, 36.5002223673027, 36.5007878662601, 36.501096365218, 
    36.5014047391758, 36.5016617391755, 36.5017442391753, 36.5018674287584, 
    36.5021073027164, 36.5024328683409, 36.502792741257, 36.5031011131315, 
    36.5032501745897, 36.5033067995896, 36.5035124339642, 36.5035405516725, 
    36.5037694881305, 36.5037866204221, 36.5039922412552, 36.5042664266714, 
    36.5047976829206, 36.5051232412534, 36.5053694902114, 36.5054144902113, 
    36.5056544881276, 36.505791551669, 36.5060657422936, 36.5064255506264, 
    36.5069346787506, 36.5069780600005, 36.5070121141671, 36.5069272391673, 
    36.5068470547924, 36.5068464881257, 36.5067511766675, 36.5064598662513, 
    36.5063913027097, 36.506456176668, 36.5065283672929, 36.5066921787509, 
    36.5067168662509, 36.5069396787506, 36.5070424870838, 36.507076739167, 
    36.5070938662503, 36.507111048542, 36.5072309256251, 36.507505180833, 
    36.5077450527077, 36.5080021162489, 36.5082419912486, 36.5085847422897, 
    36.5087046777062, 36.5089103006225, 36.5093044256219, 36.5093791787468, 
    36.5097328672879, 36.5099727402042, 36.5101098047873, 36.5102269839538, 
    36.5102468683287, 36.5104868068701, 36.5108295537445, 36.5111722433273, 
    36.5115492391601, 36.5118295516597, 36.5121832995758, 36.5125431777002, 
    36.5128516131164, 36.5131086151993, 36.5132286141575, 36.5132286162408, 
    36.5131943026992, 36.5129715506162, 36.5127828016581, 36.5126116766584, 
    36.512423178742, 36.5123203641589, 36.5124231766587, 36.5127488068666, 
    36.5130743651994, 36.5134704266571, 36.5135884308236, 36.5140511141562, 
    36.514409991239, 36.5149828631131, 36.5155199901956, 36.5158089891535, 
    36.5157899245702, 36.5157865558202, 36.5159782381115, 36.5159763026949, 
    36.5159701172782, 36.5158675526951, 36.5156104901955, 36.5152506224877, 
    36.5147708068634, 36.5142739276975, 36.5138454912399, 36.5136549891568, 
    36.5133828006155, 36.5128516151997, 36.5124403027004, 36.5120633027009, 
    36.5117476162431, 36.5114635537436, 36.5110866141608, 36.5107953037446, 
    36.5105039891617, 36.5102811777037, 36.5101098037456, 36.5100241756208, 
    36.5098870516626, 36.509681426663, 36.50942436833, 36.5092873058302, 
    36.5091330506222, 36.5090816787472, 36.509047367289, 36.5089445516641, 
    36.508841740206, 36.508773240206, 36.5088589277059, 36.5091330527055, 
    36.5095957412465, 36.5100241735374, 36.5105553652033, 36.5108099902029, 
    36.511412177702, 36.5118063047847, 36.5121318631175, 36.5123546766588, 
    36.5125088683253, 36.5126459870751, 36.5128516151997, 36.5131600547826, 
    36.5133656776989, 36.5135713620736, 36.5136398589485, 36.5136055485319, 
    36.5136055547819, 36.5136569933235, 36.5136251787402, 36.5136227412402, 
    36.5136227391569, 36.5136741162401, 36.5138208683233, 36.5138811735314, 
    36.513991990198, 36.513970618323, 36.5138283620732, 36.5136912412401, 
    36.5137084224901, 36.5137940526982, 36.5139117401981, 36.513999740198, 
    36.5142567422809, 36.5145138047805, 36.5145651776971, 36.514599483947, 
    36.514616615197, 36.5146166131137, 36.514616618322, 36.5146166110303, 
    36.5145824297804, 36.5145138026971, 36.5143766766557, 36.5142623058225, 
    36.5141368047811, 36.5140339901979, 36.5140339901979, 36.5140853620728, 
    36.5141702974893, 36.5141630537394, 36.5142443037392, 36.5144219891556, 
    36.5146000485303, 36.5146989881135, 36.514640240197, 36.5144526756139, 
    36.5142639287392, 36.514166370406, 36.513940737073, 36.5134799245737, 
    36.5132303016575, 36.5130053006162, 36.5129974308245, 36.5129646141579, 
    36.5129441183246, 36.5136623631151, 36.5139596131147, 36.5139995537396, 
    36.5142142412393, 36.5144953026972, 36.5146596797803, 36.515270993321, 
    36.5158776797784, 36.5162974901944, 36.5163674881109, 36.5164942433191, 
    36.516741492277, 36.5169471172767, 36.5170499297765, 36.5172213047763, 
    36.5174611818592, 36.5177524933171, 36.5180781151916, 36.5183694297745, 
    36.5186435526907, 36.5188149276905, 36.5188652391487, 36.5188663641487, 
    36.5188562412321, 36.5187806776905, 36.518694986024, 36.5186778651907, 
    36.518712117274, 36.518900613107, 36.5191404881066, 36.5195003641478, 
    36.5198088651889, 36.5200861162302, 36.5201175537301, 36.5203384276881, 
    36.5205386162295, 36.5208012433124, 36.5209564297705, 36.5210597391453, 
    36.5213681787282, 36.5216081151862, 36.5217451797693, 36.5217794891442, 
    36.5219019881023, 36.521903429769, 36.5222166172686, 36.522318427685, 
    36.5224435526848, 36.5230773006005, 36.5230700526839, 36.5229678662257, 
    36.5228723037258, 36.5227709266427, 36.5226968662261, 36.5226526787262, 
    36.5227203641427, 36.5229983631007, 36.5232291131003, 36.5232784922669, 
    36.5233509328918, 36.5237968683077, 36.5243958037235, 36.5247189891397, 
    36.5248780578894, 36.5250224235141, 36.5250911776807, 36.525101614139, 
    36.5250451755975, 36.5249217422643, 36.5246455568481, 36.5244744255983, 
    36.5244304901818, 36.5244083630985, 36.52447080164, 36.5245330505983, 
    36.5245368641399, 36.5245051787233, 36.5245047401817, 36.5246409297648, 
    36.5247792422646, 36.5248853630977, 36.5249640505976, 36.5251182401807, 
    36.5251328630973, 36.5253861141386, 36.5257298037214, 36.5261780537207, 
    36.5264912401786, 36.5266639912199, 36.5268001787197, 36.5273306808023, 
    36.5277500537183, 36.5280647412178, 36.5283274880924, 36.528604869342, 
    36.5287862422583, 36.5289008641332, 36.5289018641332, 36.5286488651752, 
    36.5288549891332, 36.5289219901748, 36.5289041151748, 36.5288194255916, 
    36.528582238092, 36.5284121808006, 36.5283188047591, 36.5283173662174, 
    36.5283119870508, 36.528342242259, 36.5284586724672, 36.5286604974668, 
    36.5288336787166, 36.5289026766332, 36.5289627391331, 36.5290498651746, 
    36.5290609307996, 36.5290632380912, 36.5291340547578, 36.5293719287158, 
    36.5295073672572, 36.5295475505905, 36.5295845537154, 36.5294979255905, 
    36.5293609912158, 36.5293623641325, 36.5294583672573, 36.5296777380903, 
    36.5300211766314, 36.5304029297558, 36.5306419891305, 36.5308818672551, 
    36.5311322401714, 36.5312299943379, 36.5316690526705, 36.5321542995447, 
    36.5324050526694, 36.532626490169, 36.5328186182937, 36.5331201766266, 
    36.5332885537097, 36.5336073026675, 36.5339417412087, 36.5341428037083, 
    36.5342395537082, 36.5342603651665, 36.5342543630832, 36.5343191766248, 
    36.5345053641245, 36.5347660526657, 36.5349276776655, 36.5350620526652, 
    36.5352240505817, 36.5354153651647, 36.4470129278019, 36.4471104278018, 
    36.4473000569682, 36.4476439288426, 36.4480187434253, 36.4483820538414, 
    36.4486769277993, 36.448883737174, 36.4486303611328, 36.4482023642584, 
    36.4479865528004, 36.4477123663425, 36.4476950528008, 36.447403928843, 
    36.44718117676, 36.4469926757186, 36.4467527392607, 36.4465814278026, 
    36.4465641757193, 36.446547117386, 36.4466156798859, 36.4468069903023, 
    36.4468384257189, 36.4470440507185, 36.4470440528019, 36.4468555475938, 
    36.4466793038441, 36.4466088642609, 36.4465970538442, 36.4468328642606, 
    36.4473851142597, 36.4481968028001, 36.4488510517574, 36.44931367884, 
    36.4498592434225, 36.4502381767552, 36.4507498017545, 36.4511166798789, 
    36.451244175712, 36.4512558027953, 36.4512260559204, 36.4512833642536, 
    36.4513109277952, 36.4513281184202, 36.4514137361284, 36.451670801753, 
    36.4519449902943, 36.4524590527935, 36.4527846809179, 36.4530074246676, 
    36.4533159277921, 36.4536071777917, 36.4538813632079, 36.4543093673739, 
    36.454517797582, 36.454902486123, 36.4550478632061, 36.4552146132058, 
    36.4553274913307, 36.4554096132056, 36.4553169277891, 36.4553039288307, 
    36.4553702444556, 36.4553703017473, 36.4555987444553, 36.4559032996631, 
    36.4564003017457, 36.4564378621623, 36.4566916777869, 36.457051553828, 
    36.4573429267442, 36.4573942413275, 36.457239990286, 36.4569486798698, 
    36.4567430527868, 36.4565256788288, 36.4565419267454, 36.4566418048703, 
    36.4568026757034, 36.4569311767449, 36.4570933027863, 36.4571321132029, 
    36.4573990538275, 36.4575754277855, 36.4576381788271, 36.4576513048688, 
    36.4576855548687, 36.4576098642438, 36.4575998673688, 36.4575869892439, 
    36.4573771142442, 36.4570343048697, 36.4566231111203, 36.4563832382041, 
    36.4561947402877, 36.4560949882045, 36.4560062392463, 36.4557321152884, 
    36.4553550548723, 36.4549267413313, 36.4546702413317, 36.4545124902903, 
    36.4544836777903, 36.4544824892487, 36.4545164267486, 36.454477178832, 
    36.4544982434153, 36.454481116332, 36.4545668038319, 36.4546010517485, 
    36.4546010538318, 36.4545315507069, 36.4544372434154, 36.4544870527903, 
    36.45469724029, 36.4548455517481, 36.454891426748, 36.455135616331, 
    36.4554904913304, 36.4555044871638, 36.4562008069543, 36.4564929298705, 
    36.456617490287, 36.4567655517451, 36.4569581152865, 36.4571034298696, 
    36.4571391725779, 36.4571306767446, 36.4571111767446, 36.4570032402864, 
    36.45686149237, 36.4565278017455, 36.4564049309124, 36.4562896184125, 
    36.4562441746626, 36.4560028642463, 36.4556834892468, 36.4554602402888, 
    36.4552378048725, 36.455112363206, 36.4550389882061, 36.4549718652896, 
    36.4548143038315, 36.4545919361235, 36.4543200517489, 36.4542579288324, 
    36.4539883642494, 36.4536404871666, 36.453182366334, 36.4528526163346, 
    36.452759743418, 36.4525706777933, 36.4523969892519, 36.4523836767519, 
    36.4524527382101, 36.4526813017515, 36.4526914330015, 36.4527801788346, 
    36.4529749902927, 36.4531228048758, 36.4531267382091, 36.4531283017508, 
    36.4532596757089, 36.4534546142502, 36.4537521163331, 36.4537929902914, 
    36.4538193048747, 36.4539872392494, 36.4542785538323, 36.4544842996654, 
    36.4545683684152, 36.454714680915, 36.4547101788316, 36.4547015548733, 
    36.4547363007066, 36.4547614298733, 36.4548346777898, 36.4550445548728, 
    36.4551426142476, 36.4552403027892, 36.4553852423722, 36.4557053673718, 
    36.4558448652882, 36.455980927788, 36.4560101767463, 36.456027802788, 
    36.4560933027878, 36.4561553059127, 36.4562376777876, 36.4562240527876, 
    36.4561951819543, 36.456197554871, 36.4562654871626, 36.456171114246, 
    36.4559802382047, 36.4557259257051, 36.4555513694553, 36.4550569267478, 
    36.454658362165, 36.4543076777906, 36.4540370538327, 36.4539442402912, 
    36.4536866777916, 36.4535584902918, 36.4534779288335, 36.4534121142503, 
    36.4534229330003, 36.4534563673753, 36.4533791194587, 36.4531270548758, 
    36.4528719288345, 36.4518499882111, 36.4509089246709, 36.4507026173795, 
    36.4505608632131, 36.4503224892551, 36.4501842392553, 36.4501456777971, 
    36.4496658652978, 36.4496223038395, 36.4495270538397, 36.4493060548817, 
    36.4492744267567, 36.4492648673818, 36.4492046798819, 36.4490831777987, 
    36.448894743424, 36.448671991341, 36.4486377465494, 36.4487748017575, 
    36.4489633059239, 36.4490416777988, 36.4492203652985, 36.4494431194648, 
    36.4495288048814, 36.449528802798, 36.4495174913397, 36.4494946163397, 
    36.4494088652982, 36.4494773663397, 36.4496144902979, 36.4497344298811, 
    36.4500599902972, 36.4504753652965, 36.4506644892546, 36.4510021142541, 
    36.451228300712, 36.4517432423779, 36.4521124923774, 36.4525130527934, 
    36.4528976777928, 36.4529574257094, 36.4531388642508, 36.4533019934171, 
    36.4532871777922, 36.4532723652922, 36.4532117402923, 36.4532309277923, 
    36.4534244892503, 36.4536208027916, 36.4537126163332, 36.454239864249, 
    36.4542728038323, 36.4539711757078, 36.4535581809168, 36.4530641757092, 
    36.4529056777928, 36.4527648038347, 36.4522498017521, 36.4519463017526, 
    36.4513398038369, 36.4512897402953, 36.4511053007122, 36.4507797402961, 
    36.4505398017548, 36.4505055538382, 36.4504972382132, 36.4504553027966, 
    36.4504099288383, 36.4502009288386, 36.4501903642553, 36.4502249892553, 
    36.4503605517551, 36.4504352444633, 36.4505723663381, 36.450627675713, 
    36.4506678642546, 36.4507209288378, 36.4507759892544, 36.4508256767543, 
    36.4508602361293, 36.4508676777959, 36.450835552796, 36.4507266788378, 
    36.4506316767547, 36.4504319923799, 36.4502313642553, 36.4498029892559, 
    36.4494259871732, 36.4489290548823, 36.4485863048828, 36.4483293080082, 
    36.4480551153003, 36.4480473028003, 36.4479699309255, 36.4475106153012, 
    36.4472399267599, 36.4471846132183, 36.446952612177, 36.4468100507189, 
    36.4467017340524, 36.4466499267608, 36.446547117386, 36.4464100528029, 
    36.4462215590531, 36.4459286153036, 36.4457417434289, 36.445296176763, 
    36.4451419882215, 36.4450734278049, 36.4449706194717, 36.4448335528053, 
    36.4446793059305, 36.4446793017639, 36.4447135538472, 36.4450391757217, 
    36.4452619913463, 36.4453051153046, 36.4453657403045, 36.4452882392629, 
    36.4452765538463, 36.4451623673881, 36.4449753017634, 36.4446758017639, 
    36.4441384944731, 36.4435204278074, 36.4429295517666, 36.4429169903083, 
    36.4425347382256, 36.4423076798926, 36.4418176142683, 36.4413549288524, 
    36.4411664298943, 36.4411835548943, 36.4415776778104, 36.4418861215599, 
    36.4419834288514, 36.4421599923928, 36.4422106153094, 36.4421181142679, 
    36.4420089913514, 36.4419976163514, 36.4418734934349, 36.4416386173936, 
    36.4415953048937, 36.4415779267687, 36.4417106778101, 36.4420168590597, 
    36.4423316778092, 36.4427258028086, 36.4430513632248, 36.4433941173909, 
    36.4438224944735, 36.4441138007231, 36.4442755548895, 36.4443926163477, 
    36.4445541767641, 36.444588114264, 36.4444617434309, 36.4444573028059, 
    36.444383365306, 36.4444964288475, 36.4447851163471, 36.4450900528049, 
    36.4453638038461, 36.4454949871793, 36.4455343028042, 36.4453308028046, 
    36.4448866757219, 36.4444437403059, 36.4441596142647, 36.4438212413485, 
    36.4436049319739, 36.4431914882245, 36.4425536788505, 36.4422875517676, 
    36.4419789278097, 36.4414058653106, 36.4410580517695, 36.4410454892695, 
    36.4409982330196, 36.4410546767695, 36.4411336788527, 36.4408847413531, 
    36.4408431173948, 36.4405869288536, 36.4403457996873, 36.4401500496876, 
    36.4399541736462, 36.4397281788549, 36.4393514882305, 36.4388844246895, 
    36.4384246153153, 36.4381612413573, 36.4376941778164, 36.4374229892751, 
    36.4370764309423, 36.4368138653177, 36.4364888632349, 36.4362628611519, 
    36.4361724278187, 36.4360669892773, 36.4359163017775, 36.4356300538612, 
    36.4351931778203, 36.4348164319875, 36.4344247413632, 36.4339274924056, 
    36.4335358017812, 36.433249491365, 36.432767365324, 36.4323907392829, 
    36.4319989934502, 36.4316826132424, 36.4313812413678, 36.4309443059519, 
    36.4305680507441, 36.4305073663692, 36.4299198038701, 36.4295129892874, 
    36.4292568028295, 36.4290760497047, 36.4289103674134, 36.4285789288722, 
    36.4280214278314, 36.4275694267905, 36.427207801791, 36.4269215528331, 
    36.426605117417, 36.4263942382506, 36.426153116376, 36.4258907403347, 
    36.4258668653347, 36.4256107455435, 36.4253094257523, 36.4250382392944, 
    36.4247971778364, 36.4246163632533, 36.4243753017954, 36.4241794247123, 
    36.4240588622126, 36.4240433653376, 36.4240287382543, 36.4240136726293, 
    36.4239233028377, 36.423742490338, 36.4234713028385, 36.4230042361725, 
    36.4224467434651, 36.4220372445074, 36.4217687382578, 36.4212866768002, 
    36.4209099882591, 36.4206063028429, 36.4205031757597, 36.4200059924272, 
    36.4197649288859, 36.4195690549279, 36.4193883018031, 36.4187855518041, 
    36.4184541153463, 36.4176857455558, 36.4171131799317, 36.4165858632658, 
    36.4165401778492, 36.416254364308, 36.4159379872252, 36.4155462424341, 
    36.4152136153513, 36.4149888028516, 36.4145217393107, 36.4141149268114, 
    36.4139415497282, 36.4139311768116, 36.4137126174369, 36.4133015518126, 
    36.4132502403543, 36.4132280518127, 36.4131730538961, 36.4130813674379, 
    36.4129990528547, 36.41285036223, 36.4125500528554, 36.4122146132726, 
    36.4120699913979, 36.411981738273, 36.4116876778568, 36.4113863674406, 
    36.4111151778577, 36.410859052858, 36.4105432414002, 36.4104070518171, 
    36.4102563643173, 36.4100755518176, 36.4099098039012, 36.409774239318, 
    36.4097139934848, 36.40962355286, 36.4095030507768, 36.4093523664021, 
    36.4092619914022, 36.4092921747355, 36.4094879851518, 36.4097215539015, 
    36.4097441122348, 36.4100755549426, 36.4103316778588, 36.4105727414001, 
    36.4107836747332, 36.4109343663996, 36.4110247403578, 36.4111453018159, 
    36.4113411778573, 36.4114617372321, 36.4115671768153, 36.4117479278567, 
    36.4121999257727, 36.4125464226471, 36.4126519320219, 36.4126519320219, 
    36.4125467413971, 36.4125332372304, 36.4125393695221, 36.4133766768124, 
    36.4135423663955, 36.4135875538955, 36.4134369288957, 36.4131958643127, 
    36.4129999882714, 36.4128643653549, 36.4128279268133, 36.4127890486884, 
    36.4126014903553, 36.4125630549387, 36.412404801814, 36.4123801778557, 
    36.4124191163973, 36.4126806132719, 36.413269116396, 36.4143290528527, 
    36.4153123653512, 36.4165758622242, 36.4170784288901, 36.4171583674316, 
    36.4172428018065, 36.417354243473, 36.4175350538894, 36.4176404913892, 
    36.4176857382641, 36.4176857403475, 36.4176103643059, 36.4174144872229, 
    36.4172392403481, 36.4171583643066, 36.4169624903486, 36.4168570497237, 
    36.4168570528487, 36.4169624903486, 36.4171884903482, 36.4176254278476, 
    36.4178212997222, 36.4178966143054, 36.4180322424302, 36.4182431799299, 
    36.4184842455546, 36.4186601143043, 36.4186650497209, 36.4186806143042, 
    36.4187379226375, 36.4187554299291, 36.4186801205543, 36.4184541184712, 
    36.41820886743, 36.4180924903468, 36.4176857382641, 36.4173843601396, 
    36.4171433028483, 36.417113175765, 36.4171734268066, 36.4172789278481, 
    36.417339174723, 36.4173966778479, 36.4173591163896, 36.4173948695146, 
    36.4172149903482, 36.4174366747228, 36.417723303889, 36.4178824913888, 
    36.4180267382636, 36.4186326163876, 36.419253802845, 36.4196822393027, 
    36.4199523070106, 36.4203659893016, 36.4205031809681, 36.4205031757597, 
    36.4205031788848, 36.4204881122181, 36.4204881195097, 36.4206839882594, 
    36.4210455549256, 36.4213167393002, 36.4215578632581, 36.421648238258, 
    36.4216783663829, 36.4216181153413, 36.4214975486748, 36.4214796132582, 
    36.4214638028416, 36.4213664913834, 36.4215083611749, 36.421665432008, 
    36.4217102424245, 36.4218518642993, 36.421884427841, 36.4219329267992, 
    36.4221109924239, 36.4223918059652, 36.422901113256, 36.423378048672, 
    36.4238082413796, 36.4241430486708, 36.4243982361704, 36.4244765528369, 
    36.4244583663786, 36.4245514257535, 36.4246925549199, 36.4246911788782, 
    36.4247067413782, 36.4247669882531, 36.4247434278365, 36.4246615528366, 
    36.4245108653369, 36.4244957986702, 36.42461636117, 36.4247218017949, 
    36.4248272965864, 36.4249779267944, 36.4253094278356, 36.4255242392936, 
    36.4255546153352, 36.4259056809597, 36.4261600549176, 36.4262544309591, 
    36.4262516747091, 36.4260727361678, 36.4257178663767, 36.4249634267945, 
    36.4247566153365, 36.4245492434618, 36.4245396205452, 36.4242456153373, 
    36.4240059892959, 36.4237819299213, 36.4236052392966, 36.4233163653387, 
    36.4231074267973, 36.4229460528393, 36.4229609892976, 36.4231670538806, 
    36.4231978028389, 36.4230997403391, 36.4230663632558, 36.4230968080474, 
    36.423335742422, 36.4234133632552, 36.4236022392966, 36.4237095517964, 
    36.4237870538797, 36.4238968090878, 36.4237039267965, 36.4233995528386, 
    36.4233272434637, 36.4230940549224, 36.4230291122142, 36.4230273632558, 
    36.4230739257558, 36.4232643007555, 36.4235318028384, 36.4238753663795, 
    36.424198741379, 36.4245014267952, 36.4247868642947, 36.4249260580445, 
    36.4250671195027, 36.4250903038776, 36.4254476820021, 36.4257339278349, 
    36.4261487392927, 36.42676980075, 36.4271470517911, 36.4275240528322, 
    36.427401053874, 36.427415928874, 36.4277648038735, 36.427808929915, 
    36.4280986142896, 36.4281928038728, 36.428316487206, 36.428285618456, 
    36.4282624913727, 36.4279309924149, 36.4277954257484, 36.4279159236649, 
    36.4279755507482, 36.4280364278314, 36.4280364257481, 36.4280364257481, 
    36.4279761819981, 36.4279761809565, 36.4279761767898, 36.4280063684564, 
    36.4281721194978, 36.4283227372059, 36.4283696174142, 36.4284996132473, 
    36.4289706767883, 36.4289876153299, 36.4291440538713, 36.4294479267875, 
    36.4295589299123, 36.4295724861623, 36.4297917382453, 36.4298403642869, 
    36.4298688684535, 36.4300253028283, 36.4304994913692, 36.4307199299105, 
    36.430895427827, 36.4310697319933, 36.4311950528265, 36.4314804882427, 
    36.4317649892839, 36.4319057361587, 36.4320324288668, 36.4320471726168, 
    36.4319166153253, 36.4319308049087, 36.431931366367, 36.431947241367, 
    36.4321643007416, 36.4322012403249, 36.4323456799081, 36.4327748642824, 
    36.4330775517819, 36.433426177823, 36.433435302823, 36.433673801781, 
    36.4338672371973, 36.4341233642803, 36.4342136132385, 36.4343493621966, 
    36.4346054871962, 36.4348179278209, 36.4348616194874, 36.4350725507371, 
    36.4353286757367, 36.4354341767782, 36.4355698028197, 36.4357656174027, 
    36.4360519299022, 36.4362025507353, 36.4362326778187, 36.4360971121939, 
    36.4357958028193, 36.4355315496948, 36.4352432996952, 36.4350485507372, 
    36.4350126163622, 36.4349499257373, 36.434945551779, 36.434910929904, 
    36.4350110507372, 36.4352621819868, 36.4351151142787, 36.4350934278204, 
    36.4350584955288, 36.4349932382373, 36.4349439871957, 36.4348971778207, 
    36.4348769288624, 36.434715802821, 36.4343480507383, 36.4342271174051, 
    36.4338203059474, 36.4334844892813, 36.4331806757401, 36.4330836767819, 
    36.4330498038653, 36.4330021153237, 36.4329992371987, 36.4329919278237, 
    36.4329082392821, 36.4328863049072, 36.4325983007409, 36.4324851153245, 
    36.4324059236579, 36.4323883059496, 36.4322924288664, 36.4322793674081, 
    36.4320830517834, 36.4324080517829, 36.4327169267825, 36.4329899215737, 
    36.4332509882399, 36.4334933674062, 36.4335436153228, 36.4338286788641, 
    36.4339525517805, 36.4339783007388, 36.4340146767804, 36.4340369861554, 
    36.434082490322, 36.4341274934469, 36.4343376184466, 36.4344163653215, 
    36.4343826184465, 36.4343092413633, 36.4342691778217, 36.4341404965719, 
    36.4340431132387, 36.4339831778221, 36.4339805507388, 36.4339134882389, 
    36.4338233049057, 36.4337568028225, 36.4342046142801, 36.43430305178, 
    36.4342540528218, 36.4343391757383, 36.434504863238, 36.4346486153211, 
    36.4349611163623, 36.4351774924036, 36.4353549892784, 36.4356946153195, 
    36.4358951153192, 36.4357587382361, 36.435566617403, 36.435604673653, 
    36.4358772403192, 36.4363247371935, 36.4364460528183, 36.4364859913599, 
    36.4364562371933, 36.4365689924015, 36.4363815549017, 36.4361094871938, 
    36.4358061778193, 36.435581614278, 36.4354211788616, 36.4352455496952, 
    36.4350374257372, 36.4347487392793, 36.4345548049046, 36.434516681988, 
    36.4344201746965, 36.4342592403217, 36.4342093049052, 36.4342048663635, 
    36.4341914267802, 36.43430055178, 36.43428310803, 36.4342329299051, 
    36.4340922392803, 36.4340903632386, 36.433898613239, 36.4333663069898, 
    36.4330683621986, 36.432981739282, 36.4327959892823, 36.4324907382411, 
    36.4322664299082, 36.4319138049087, 36.4315438632426, 36.431504927826, 
    36.4312199267848, 36.4311797361598, 36.4312263049098, 36.4313623674096, 
    36.4315550486593, 36.4317624892839, 36.4318462392838, 36.431961738242, 
    36.4321829924083, 36.4324721142828, 36.4325622455327, 36.4330054903237, 
    36.4333398642815, 36.4335553017812, 36.4335793632395, 36.4337333674059, 
    36.4338829246973, 36.4340254913637, 36.4343606726133, 36.4347082424044, 
    36.4353028674034, 36.4355587392781, 36.4358710538609, 36.436861989276, 
    36.4375877371916, 36.4382399236489, 36.4386704882315, 36.4387501767731, 
    36.4389444913561, 36.4390273048976, 36.4391073642725, 36.4391254923975, 
    36.4393186726055, 36.4394173663554, 36.4395134288552, 36.4397203048966, 
    36.4399749246879, 36.4403588028122, 36.4406951173951, 36.4408009913532, 
    36.4408555538532, 36.4411239913528, 36.4415163028104, 36.4422938684343, 
    36.4427257392669, 36.443062052808, 36.4432216778078, 36.4433807403076, 
    36.4435228653073, 36.4439239903067, 36.4441813048896, 36.4444075507226, 
    36.4447937392637, 36.4450832392632, 36.4451471798882, 36.4455469913459, 
    36.4460283673868, 36.4463290507197, 36.4464730538444, 36.4465543653026, 
    36.4465689903026, 36.4465725517609, 36.4467276767607, 36.4470129278019 ;

 geometry_container = _ ;

 node_count = 1678, 950 ;

 crs = _ ;
}
