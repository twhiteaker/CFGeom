netcdf multiline_vlen {
types:
  double(*) node_VLType ;
  int(*) part_node_VLType ;
dimensions:
	instance = 2 ;
variables:
	int geometry_container ;
		geometry_container:geometry_type = "line" ;
		geometry_container:node_coordinates = "x y" ;
		geometry_container:part_node_count = "part_node_count" ;
	node_VLType x(instance) ;
		x:axis = "X" ;
	node_VLType y(instance) ;
		y:axis = "Y" ;
	part_node_VLType part_node_count(instance) ;
		part_node_count:long_name = "count of nodes in each geometry part" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 geometry_container = _ ;

 x = {3, 1, 4}, {1, 2, 4, 3} ;

 y = {1, 3, 4}, {2, 4, 3, 2} ;

 part_node_count = {3}, {2, 2} ;
}
