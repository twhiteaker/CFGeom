netcdf file\:/C\:/Temp/dsg/nwm_bullcreek {
  dimensions:
    time = 1;
    station = 20;
  variables:
    int time(time);
      time:units = "seconds since 2016-05-26 06:00 UTC";
      time:long_name = "valid output time";

    int station_id(station);
      station_id:long_name = "Station id";

    double streamflow(station);
      streamflow:long_name = "River Flow";
      streamflow:units = "meter^3 / sec";

  // global attributes:
  :Conventions = "Unidata Observation Dataset v1.0";
  :cdm_datatype = "Station";
  :model_initialization_time = "2016-05-26_06:00:00";
  :station_dimension = "station";
  :missing_value = -8.9999998E15f;
  :stream_order_output = 1;
  :model_output_valid_time = "2016-05-27_00:00:00";
 data:
time =
  {21600}
station_id =
  {5781157, 5781193, 5781183, 5781189, 5781173, 5781133, 5781163, 5781131, 5781141, 5781171, 5781159, 5781129, 5781139, 5781149, 5781185, 5781187, 5781145, 5781781, 5781191, 5781811}
streamflow =
  {0.25217628479003906, 0.0201607346534729, 0.03469820320606232, 0.06074899435043335, 0.08355419337749481, 0.3565440773963928, 0.1054951474070549, 0.07029025256633759, 0.21661187708377838, 0.03520715981721878, 0.03696829080581665, 0.10193829983472824, 0.12274756282567978, 0.37541332840919495, 0.6298931241035461, 0.7174544930458069, 1.1098110675811768, 1.1597568988800049, 1.3793467283248901, -1.999399951158054E-11}
}
