netcdf point_z_vlen {
dimensions:
	instance = 2 ;
variables:
	int geometry_container ;
		geometry_container:geometry_type = "point" ;
		geometry_container:node_coordinates = "x y z" ;
	double x(instance) ;
		x:axis = "X" ;
	double y(instance) ;
		y:axis = "Y" ;
	double z(instance) ;
		z:axis = "Z" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 geometry_container = _ ;

 x = 1, 2 ;

 y = 1, 3 ;

 z = NaN, 50 ;
}
