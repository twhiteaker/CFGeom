netcdf line_cra {
dimensions:
	instance = 2 ;
	node = 5 ;
variables:
	int geometry_container ;
		geometry_container:geometry_type = "line" ;
		geometry_container:node_coordinates = "x y" ;
		geometry_container:node_count = "node_count" ;
	double x(node) ;
		x:axis = "X" ;
	double y(node) ;
		y:axis = "Y" ;
	int node_count(instance) ;
		node_count:long_name = "count of coordinates in each instance geometry" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 geometry_container = _ ;

 x = 3, 1, 4, 7, 8 ;

 y = 1, 3, 4, 9, 10 ;

 node_count = 3, 2 ;
}
