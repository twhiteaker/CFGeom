netcdf polygon_hole_vlen {
types:
  double(*) node_VLType ;
  int(*) part_node_VLType ;
dimensions:
	instance = 2 ;
variables:
	int geometry_container ;
		geometry_container:geometry_type = "polygon" ;
		geometry_container:node_coordinates = "x y" ;
		geometry_container:part_node_count = "part_node_count" ;
		geometry_container:interior_ring = "interior_ring" ;
	node_VLType x(instance) ;
		x:axis = "X" ;
	node_VLType y(instance) ;
		y:axis = "Y" ;
	part_node_VLType part_node_count(instance) ;
		part_node_count:long_name = "count of nodes in each geometry part" ;
	part_node_VLType interior_ring(instance) ;
		interior_ring:long_name = "type of each polygon geometry part" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 geometry_container = _ ;

 x = {10, 5, 0, 1, 5, 9}, {20, 15, 11, 15} ;

 y = {0, 5, 0, 1, 4, 1}, {20, 25, 20, 15} ;

 part_node_count = {3, 3}, {4} ;

 interior_ring = {0, 1}, {0} ;
}
