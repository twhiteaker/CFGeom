netcdf bull_creek_with_geom_CRA {
dimensions:
	time = 15 ;
	comid = 20 ;
	flowlines_node = 515 ;
	flowlines_GNIS_NAME_strlen = 15 ;
	catchments_node = 4275 ;
	catchments_part = 21 ;
variables:
	int time(time) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 2016-11-07 20:00 UTC" ;
	int comid(comid) ;
		comid:cf_role = "timeseries_id" ;
	double lat(comid) ;
		lat:long_name = "Latitude of upstream end of river segment" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
	double lon(comid) ;
		lon:long_name = "Longitude of upstream end of river segment" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
	float streamflow(time, comid) ;
		streamflow:long_name = "River Flow" ;
		streamflow:units = "meter^3 / sec" ;
		streamflow:missing_value = -9.e+015f ;
		streamflow:coordinates = "time lat lon" ;
		streamflow:grid_mapping = "crs" ;
		streamflow:geometry = "flowlines_geometry_container" ;
	int crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;
	int flowlines_geometry_container ;
		flowlines_geometry_container:geometry_type = "line" ;
		flowlines_geometry_container:node_coordinates = "flowlines_x flowlines_y flowlines_z" ;
		flowlines_geometry_container:node_count = "flowlines_node_count" ;
	double flowlines_x(flowlines_node) ;
		flowlines_x:axis = "X" ;
	double flowlines_y(flowlines_node) ;
		flowlines_y:axis = "Y" ;
	double flowlines_z(flowlines_node) ;
		flowlines_z:axis = "Z" ;
	int flowlines_node_count(comid) ;
		flowlines_node_count:long_name = "count of coordinates in each instance geometry" ;
	char flowlines_GNIS_NAME(comid, flowlines_GNIS_NAME_strlen) ;
	int catchments_geometry_container ;
		catchments_geometry_container:geometry_type = "polygon" ;
		catchments_geometry_container:node_coordinates = "catchments_x catchments_y" ;
		catchments_geometry_container:node_count = "catchments_node_count" ;
		catchments_geometry_container:part_node_count = "catchments_part_node_count" ;
	double catchments_x(catchments_node) ;
		catchments_x:axis = "X" ;
	double catchments_y(catchments_node) ;
		catchments_y:axis = "Y" ;
	int catchments_node_count(comid) ;
		catchments_node_count:long_name = "count of coordinates in each instance geometry" ;
	int catchments_part_node_count(catchments_part) ;
		catchments_part_node_count:long_name = "count of nodes in each geometry part" ;
	double catchments_AreaSqKM(comid) ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:featureType = "timeSeries" ;
data:

 time = 0, 3600, 7200, 10800, 14400, 18000, 21600, 25200, 28800, 32400, 
    36000, 39600, 43200, 46800, 50400 ;

 comid = 5781157, 5781193, 5781183, 5781189, 5781173, 5781133, 5781163, 
    5781131, 5781141, 5781171, 5781159, 5781129, 5781139, 5781149, 5781185, 
    5781187, 5781145, 5781781, 5781191, 5781811 ;

 lat = 30.394875219, 30.35987842, 30.382667486, 30.37520702, 30.390782686, 
    30.419268819, 30.418718086, 30.419385019, 30.412698819, 30.421760686, 
    30.419293419, 30.449735086, 30.413898419, 30.402990419, 30.395374286, 
    30.385456486, 30.411992219, 30.411970019, 30.37150722, 30.35836542 ;

 lon = -97.839571625, -97.788739225, -97.770506225, -97.784337692, 
    -97.773616625, -97.807644692, -97.806455225, -97.810685625, 
    -97.822483092, -97.766602225, -97.776045225, -97.826984892, 
    -97.845698425, -97.848716292, -97.825136825, -97.841002625, 
    -97.832187625, -97.834487892, -97.804296025, -97.788106425 ;

 streamflow =
  0.01282661, 0.4214232, 0.6132626, 0.3697329, 0.2777951, 0.07792676, 
    0.2128945, 0.02207282, 0.02037233, 0.2944577, 0.05495298, 0.05580963, 
    0.001649335, 0.006848401, 0.01060254, 0.02235815, 0.007151061, 
    0.006909644, 0.04669686, -9e+015,
  0.0128412, 0.30901, 0.2857758, 0.2768533, 0.1787811, 0.07953472, 0.1490608, 
    0.02223668, 0.02054201, 0.1020646, 0.02873886, 0.05726831, 0.001643664, 
    0.007000346, 0.0107078, 0.005730267, 0.007306212, 0.007061725, 
    0.03053636, -9e+015,
  0.01294264, 0.2950936, 0.2652008, 0.2710669, 0.1718954, 0.07931047, 
    0.1389588, 0.02236207, 0.02085562, 0.09134504, 0.03269129, 0.0569133, 
    0.001459687, 0.007241051, 0.01085213, 0.008282697, 0.007551769, 
    0.007302842, 0.02308411, -9e+015,
  0.01302564, 0.2963086, 0.2631511, 0.2726015, 0.1623622, 0.0797341, 
    0.1433699, 0.02247054, 0.02096333, 0.09949419, 0.01842695, 0.05722875, 
    0.001460453, 0.00726573, 0.01092073, 0.008298121, 0.007576539, 
    0.007327508, 0.02320509, -9e+015,
  0.01310898, 0.3007611, 0.2649506, 0.276682, 0.1634004, 0.08016156, 
    0.1442623, 0.02257986, 0.02107178, 0.1000877, 0.01851827, 0.0575469, 
    0.001461336, 0.007290781, 0.01098949, 0.008349704, 0.007601709, 
    0.00735255, 0.02335536, -9e+015,
  0.01319266, 0.3042439, 0.2666953, 0.2799444, 0.1643, 0.08059214, 0.145032, 
    0.02268989, 0.02118085, 0.1009216, 0.01864383, 0.05786745, 0.0014623, 
    0.007316067, 0.0110585, 0.008401643, 0.007627148, 0.007377835, 
    0.02350691, -9e+015,
  0.01327646, 0.3161424, 0.272208, 0.2861931, 0.1676358, 0.08102527, 
    0.1481796, 0.0228003, 0.02129028, 0.1030719, 0.01877265, 0.05819018, 
    0.001463286, 0.007341582, 0.01150162, 0.01369355, 0.007652818, 
    0.00740335, 0.02926836, -9e+015,
  0.01336032, 0.3105679, 0.2705468, 0.2857255, 0.1662269, 0.08146068, 
    0.146677, 0.02291094, 0.02139991, 0.1027254, 0.01890479, 0.05851495, 
    0.001464299, 0.007367246, 0.01119281, 0.00850965, 0.007678639, 
    0.007429013, 0.02381739, -9e+015,
  0.01344416, 0.312577, 0.2721182, 0.2877026, 0.1669867, 0.08189801, 
    0.147381, 0.02302177, 0.0215097, 0.1036264, 0.01904018, 0.05884145, 
    0.001465337, 0.007393077, 0.01126608, 0.0085588, 0.007704631, 
    0.007454843, 0.02396684, -9e+015,
  0.01352791, 0.3150007, 0.2739817, 0.2899553, 0.1679883, 0.08233685, 
    0.1481747, 0.02313267, 0.02161955, 0.1044905, 0.01917857, 0.0591694, 
    0.001466401, 0.007419034, 0.01133522, 0.008611545, 0.00773075, 0.0074808, 
    0.02412144, -9e+015,
  0.01361153, 0.4016319, 0.3468528, 0.3696412, 0.1715118, 0.08277698, 
    0.1489779, 0.02324354, 0.02172934, 0.163293, 0.01931971, 0.05949866, 
    0.001467487, 0.00744508, 0.01141543, 0.008664394, 0.007756962, 
    0.007506847, 0.02971038, -9e+015,
  0.8212371, 12.75619, 1.100087, 0.9671487, 1.255758, 6.353597, 1.987978, 
    6.037886, 5.872139, 0.2936869, 0.08297366, 1.294393, 1.352076, 9.051786, 
    2.018898, 16.95288, 9.056293, 9.399705, 14.4407, -9e+015,
  2.142261, 14.99611, 5.313879, 3.025236, 9.933393, 16.23151, 11.75364, 
    11.43945, 8.575498, 0.2237048, 0.05611701, 5.09092, 2.952026, 3.791275, 
    4.098896, 7.154664, 5.000048, 4.010376, 12.19778, -9e+015,
  3.098789, 19.56161, 14.09752, 13.04749, 14.25079, 12.50853, 14.09196, 
    8.301886, 5.8725, 0.09821253, 0.03662128, 4.073664, 2.357652, 2.158805, 
    3.0272, 2.892411, 2.463751, 2.223096, 6.78826, -9e+015,
  2.43078, 17.1487, 14.61003, 14.3829, 14.76154, 14.10111, 14.82771, 
    6.887359, 4.316349, 0.1081519, 0.02483639, 7.233815, 2.537459, 0.9709879, 
    1.404317, 0.6012301, 1.328571, 1.032546, 2.658216, -9e+015 ;

 crs = _ ;

 flowlines_geometry_container = _ ;

 flowlines_x = -97.839571625, -97.8381966919999, -97.837403492, 
    -97.8355788919999, -97.834283092, -97.8332516249999, -97.832934225, 
    -97.8325106249999, -97.8321928249999, -97.8319812249999, -97.831531492, 
    -97.829389492, -97.827168092, -97.826533292, -97.8261362919999, 
    -97.824813825, -97.824152425, -97.823649625, -97.823411492, 
    -97.823066625, -97.823065825, -97.822483625, -97.8223776249999, 
    -97.822403825, -97.822483092, -97.788739225, -97.7884224919999, 
    -97.7882118919999, -97.788106425, -97.770506225, -97.770823692, 
    -97.7720140919999, -97.773363492, -97.773893025, -97.774238092, 
    -97.774476292, -97.775005425, -97.7754020249999, -97.7761422249999, 
    -97.776380025, -97.7781500249999, -97.7798674919999, -97.7809244919999, 
    -97.781294625, -97.782140692, -97.782590292, -97.7834898249999, 
    -97.783992825, -97.784337692, -97.784337692, -97.784391892, 
    -97.784578292, -97.785399492, -97.7854528249999, -97.7857178249999, 
    -97.785639025, -97.785190625, -97.785191092, -97.785323625, 
    -97.786063825, -97.7868832249999, -97.7878080249999, -97.788046025, 
    -97.788601625, -97.788998625, -97.7893430249999, -97.789317492, 
    -97.789055092, -97.7889758919999, -97.788950025, -97.788791692, 
    -97.788739225, -97.773616625, -97.771714092, -97.771344492, 
    -97.770764092, -97.770422292, -97.7703448249999, -97.770506225, 
    -97.8076446919999, -97.807142492, -97.806693025, -97.806455225, 
    -97.806455225, -97.803150825, -97.801934425, -97.801220292, 
    -97.798575425, -97.797252892, -97.7948722249999, -97.794131692, 
    -97.7932590249999, -97.7930210919999, -97.792862692, -97.792863225, 
    -97.792969225, -97.793472292, -97.794081025, -97.794583625, 
    -97.795218625, -97.795589225, -97.795589825, -97.795457825, 
    -97.7948502249999, -97.793080225, -97.792842625, -97.792737292, 
    -97.7927118919999, -97.793189892, -97.7933494919999, -97.793351625, 
    -97.793245892, -97.792691092, -97.792056692, -97.7916336919999, 
    -97.790391025, -97.786768492, -97.785949092, -97.785579092, 
    -97.784733692, -97.783836225, -97.783809892, -97.783678025, 
    -97.782940292, -97.782518292, -97.7819636249999, -97.781435092, 
    -97.7802986249999, -97.776862092, -97.776518892, -97.776439825, 
    -97.7764138919999, -97.776705825, -97.777553492, -97.777844825, 
    -97.778797492, -97.7791946249999, -97.779247825, -97.7790894249999, 
    -97.778640092, -97.777873492, -97.775176892, -97.7748330919999, 
    -97.774145425, -97.773616625, -97.810685625, -97.810156892, 
    -97.8094694919999, -97.808491025, -97.8076446919999, -97.822483092, 
    -97.821424225, -97.820551225, -97.818699892, -97.817324625, 
    -97.814837892, -97.813727025, -97.811399825, -97.810685625, 
    -97.766602225, -97.764937292, -97.760364492, -97.760047492, 
    -97.758991425, -97.7580676919999, -97.757408025, -97.757144825, 
    -97.756909025, -97.756698292, -97.7566190919999, -97.756566492, 
    -97.756249625, -97.756171625, -97.755089025, -97.754508492, 
    -97.7542712919999, -97.754271892, -97.7545368249999, -97.754881025, 
    -97.757791625, -97.7582944919999, -97.758903692, -97.7591692249999, 
    -97.759487092, -97.761181225, -97.761974825, -97.763191292, 
    -97.763403225, -97.763457225, -97.763168892, -97.763089625, 
    -97.763064892, -97.7631710919999, -97.7638602919999, -97.765024625, 
    -97.765554225, -97.7657402249999, -97.7658206249999, -97.765715825, 
    -97.765954692, -97.7664310919999, -97.767462625, -97.768124225, 
    -97.768839892, -97.769501492, -97.7698980919999, -97.770506225, 
    -97.776045225, -97.7757812249999, -97.775069225, -97.774145092, 
    -97.773855025, -97.773696692, -97.7733282249999, -97.773090892, 
    -97.772509825, -97.772404692, -97.7723254919999, -97.772168092, 
    -97.772142625, -97.7724082249999, -97.772620225, -97.773043625, 
    -97.773520492, -97.773547625, -97.773311092, -97.773231825, 
    -97.773205692, -97.7728628249999, -97.7723348919999, -97.772150225, 
    -97.771808692, -97.7716240249999, -97.770937492, -97.770568092, 
    -97.770146692, -97.769936692, -97.7699900919999, -97.770334292, 
    -97.770889892, -97.772317825, -97.773640292, -97.7738520249999, 
    -97.7739582249999, -97.773880025, -97.773774692, -97.773695425, 
    -97.773616625, -97.826984892, -97.8255042919999, -97.8245526919999, 
    -97.823918092, -97.823548025, -97.821749692, -97.821115225, 
    -97.819423625, -97.819317892, -97.818762825, -97.818445692, 
    -97.8174150249999, -97.816912825, -97.815247625, -97.8146136249999, 
    -97.814164825, -97.814085825, -97.814086692, -97.8144320919999, 
    -97.8146968249999, -97.815622892, -97.815834625, -97.815887692, 
    -97.8157820919999, -97.8149626919999, -97.8147250919999, 
    -97.8146988249999, -97.814619425, -97.814593025, -97.814804892, 
    -97.814831692, -97.814171092, -97.814171492, -97.814648425, 
    -97.8146488249999, -97.814305425, -97.812772492, -97.8121116249999, 
    -97.810234092, -97.8095730919999, -97.809123692, -97.808542425, 
    -97.808040492, -97.8076446919999, -97.845698425, -97.844984492, 
    -97.8443762919999, -97.843450892, -97.843001425, -97.842340625, 
    -97.842049692, -97.841124225, -97.8402514919999, -97.839801892, 
    -97.839140625, -97.838637892, -97.837765092, -97.837394825, 
    -97.8368392249999, -97.8361776249999, -97.835701292, -97.8351986919999, 
    -97.834458092, -97.833611892, -97.831681825, -97.830518292, 
    -97.829804225, -97.8290106919999, -97.828111625, -97.826789425, 
    -97.825969492, -97.8255728249999, -97.824779092, -97.824197225, 
    -97.820838825, -97.820045425, -97.819516425, -97.818511692, 
    -97.817824092, -97.817242092, -97.816898425, -97.8163168249999, 
    -97.814704292, -97.813567425, -97.8125362919999, -97.811531492, 
    -97.811002692, -97.810685625, -97.8487162919999, -97.847076492, 
    -97.846944225, -97.846705825, -97.846573425, -97.846203225, 
    -97.845885825, -97.845489292, -97.844537492, -97.843770892, 
    -97.843427092, -97.842792425, -97.840941292, -97.840042092, 
    -97.839381025, -97.836736692, -97.836392825, -97.836154492, 
    -97.8359164249999, -97.8348052919999, -97.834487892, -97.825136825, 
    -97.824528825, -97.824132092, -97.8210646919999, -97.820086292, 
    -97.819001892, -97.818631625, -97.817706292, -97.816199492, 
    -97.8154330249999, -97.8147988919999, -97.8143760249999, -97.813292092, 
    -97.812393625, -97.810517025, -97.809645092, -97.809222625, 
    -97.808932425, -97.809039292, -97.808907292, -97.807691625, 
    -97.807189492, -97.8069518249999, -97.806925625, -97.807243292, 
    -97.807878225, -97.807878492, -97.807218425, -97.807060092, 
    -97.806743292, -97.8063734249999, -97.806214892, -97.805211092, 
    -97.804259825, -97.804312892, -97.8046304919999, -97.8046572919999, 
    -97.804499092, -97.803839425, -97.8038132249999, -97.803734025, 
    -97.803709225, -97.804477492, -97.804372692, -97.804400092, 
    -97.804506225, -97.804506625, -97.804295625, -97.804296025, 
    -97.841002625, -97.840447625, -97.839205292, -97.838756025, 
    -97.838306825, -97.836509625, -97.836086892, -97.835769892, 
    -97.835241692, -97.8349512249999, -97.834159292, -97.8337102249999, 
    -97.8312524249999, -97.829720025, -97.829033092, -97.828293425, 
    -97.825705092, -97.824437292, -97.823935492, -97.823512825, 
    -97.823063492, -97.821873892, -97.821212825, -97.821133425, 
    -97.820869025, -97.8204196249999, -97.8197062249999, -97.8191774919999, 
    -97.817036425, -97.814551492, -97.812965492, -97.811776292, 
    -97.8115648249999, -97.810136492, -97.8095284249999, -97.808920492, 
    -97.807519692, -97.806859225, -97.805220692, -97.8045338919999, 
    -97.804296025, -97.832187625, -97.8315530249999, -97.830838892, 
    -97.829622292, -97.829172692, -97.8278506249999, -97.8273216919999, 
    -97.826370025, -97.8252860919999, -97.824360825, -97.823673292, 
    -97.822615425, -97.822483092, -97.834487892, -97.8343838919999, 
    -97.834120892, -97.832661292, -97.832326892, -97.832187625, 
    -97.804296025, -97.8042698249999, -97.803794492, -97.8028442249999, 
    -97.8025536919999, -97.8022368919999, -97.8014186249999, 
    -97.8006262919999, -97.7999656919999, -97.799384225, -97.798088825, 
    -97.7974542919999, -97.7962386249999, -97.795921492, -97.795446225, 
    -97.7952352249999, -97.795024425, -97.7949986249999, -97.795130892, 
    -97.795421892, -97.796506025, -97.796744292, -97.7964536919999, 
    -97.794894292, -97.794524425, -97.793758425, -97.793467892, 
    -97.793203892, -97.793072425, -97.792676425, -97.791963225, 
    -97.7912234249999, -97.790219225, -97.789294092, -97.788739225, 
    -97.788106425, -97.788017692, -97.787525492, -97.785169825, 
    -97.7838350919999, -97.783535225, -97.783513292, -97.783931692, 
    -97.784793092, -97.786389292, -97.789449425, -97.790319025, 
    -97.791174892, -97.791741825 ;

 flowlines_y = 30.394875219, 30.395149819, 30.395470286, 30.3963864190001, 
    30.397211219, 30.3981274860001, 30.3985170190001, 30.399548086, 
    30.400831419, 30.401243886, 30.4016562190001, 30.4025720860001, 
    30.4036712860001, 30.4041294190001, 30.404908419, 30.4058474190001, 
    30.4066034860001, 30.407336619, 30.4078634860001, 30.4097196860001, 
    30.4109802190001, 30.411919486, 30.4122174190001, 30.412652886, 
    30.4126988190001, 30.35987842, 30.3593740860001, 30.3585258860001, 
    30.35836542, 30.3826674860001, 30.382301086, 30.38147702, 
    30.3802406200001, 30.3794618860001, 30.3781100200001, 30.377743486, 
    30.3772624860001, 30.3770796200001, 30.377011286, 30.37705742, 
    30.37795262, 30.3787100860001, 30.3789630860001, 30.378963286, 
    30.37864302, 30.378276686, 30.37738362, 30.3766276200001, 
    30.3752070200001, 30.3752070200001, 30.3738548860001, 30.3725028860001, 
    30.37041802, 30.3699368860001, 30.3692266200001, 30.3686308200001, 
    30.3677136860001, 30.36714082, 30.36688882, 30.3666372860001, 
    30.36656902, 30.3666612860001, 30.3665698200001, 30.36597442, 
    30.36528702, 30.36437062, 30.363270486, 30.3611848200001, 30.361047286, 
    30.3605662200001, 30.3602680860001, 30.35987842, 30.3907826860001, 
    30.3900248190001, 30.389612019, 30.3885802190001, 30.3868382860001, 
    30.385211086, 30.3826674860001, 30.419268819, 30.418993486, 30.418901486, 
    30.4187180860001, 30.4187180860001, 30.417547486, 30.417501019, 
    30.4176608860001, 30.418530086, 30.418896019, 30.4198570190001, 
    30.419971086, 30.4199704860001, 30.4198558190001, 30.419626486, 
    30.4190766190001, 30.4187558190001, 30.417999819, 30.417473086, 
    30.417221419, 30.416740486, 30.4163052860001, 30.4156178860001, 
    30.415319819, 30.4145860190001, 30.412843219, 30.412430419, 
    30.4118116860001, 30.410757419, 30.4084890190001, 30.4071370190001, 
    30.4049140860001, 30.4047306190001, 30.4042718860001, 30.4040652190001, 
    30.4040648860001, 30.404270286, 30.4045428860001, 30.404404819, 
    30.4042212190001, 30.4035102190001, 30.4021344860001, 30.401882286, 
    30.4016530860001, 30.3989024860001, 30.397916686, 30.397412086, 
    30.397205619, 30.396952619, 30.3966290860001, 30.396216286, 30.395964086, 
    30.395437019, 30.394474686, 30.392596219, 30.3921838860001, 
    30.3912450190001, 30.3906724190001, 30.390282819, 30.390099419, 
    30.3899844860001, 30.3899610190001, 30.390211019, 30.3903024190001, 
    30.3906456190001, 30.3907826860001, 30.4193850190001, 30.4191784860001, 
    30.4190406860001, 30.4190630190001, 30.419268819, 30.4126988190001, 
    30.4148754190001, 30.415677219, 30.416180486, 30.4167070190001, 
    30.418264219, 30.418699019, 30.419110286, 30.4193850190001, 30.421760686, 
    30.4209572190001, 30.419394686, 30.4190964860001, 30.4177892860001, 
    30.4163676860001, 30.4151752860001, 30.4143042860001, 30.4125164860001, 
    30.411851686, 30.4118058190001, 30.4115536190001, 30.4111866860001, 
    30.410201219, 30.409008419, 30.408091219, 30.4074952190001, 
    30.4070138860001, 30.406578686, 30.406235419, 30.404404619, 30.403900886, 
    30.403053619, 30.402160086, 30.4015874190001, 30.399801419, 
    30.3994354860001, 30.399092819, 30.3987722190001, 30.397832619, 
    30.3957926860001, 30.395723886, 30.394211419, 30.393890619, 
    30.3921724190001, 30.391279619, 30.390455219, 30.3896760860001, 
    30.388667819, 30.387865619, 30.387017886, 30.386537086, 30.3860566860001, 
    30.385369686, 30.3834682200001, 30.3828040860001, 30.3826898200001, 
    30.3826674860001, 30.419293419, 30.418880819, 30.4171156190001, 
    30.4157626860001, 30.4149604190001, 30.414708219, 30.4131494860001, 
    30.4125306190001, 30.4120030190001, 30.4113840860001, 30.4113154190001, 
    30.4101694190001, 30.409275619, 30.408129886, 30.407671819, 
    30.4072596190001, 30.4064348860001, 30.4057474860001, 30.4045556190001, 
    30.404509686, 30.404188886, 30.4034094190001, 30.4026984860001, 
    30.402308686, 30.400223086, 30.3999020860001, 30.3990764860001, 
    30.3984574190001, 30.3970132860001, 30.395661019, 30.3952026860001, 
    30.394721686, 30.3944014190001, 30.3940358190001, 30.3933952190001, 
    30.3931892190001, 30.3927538190001, 30.391607886, 30.3912182190001, 
    30.391172286, 30.3907826860001, 30.449735086, 30.448244819, 30.447190219, 
    30.4466628860001, 30.4464564190001, 30.4457682190001, 30.4453782860001, 
    30.4434524860001, 30.4431774190001, 30.4425584190001, 30.442031086, 
    30.4408388860001, 30.4404262190001, 30.4387752860001, 30.437720819, 
    30.436506019, 30.435818419, 30.4343516860001, 30.4321518190001, 
    30.431716486, 30.431098219, 30.430846219, 30.430525419, 30.4303190860001, 
    30.4295852860001, 30.429149819, 30.4289206190001, 30.428874819, 
    30.4286684190001, 30.428233086, 30.4276374190001, 30.4268348860001, 
    30.426216219, 30.4250476190001, 30.4244516860001, 30.4239474190001, 
    30.4226174190001, 30.4223420860001, 30.422295219, 30.422134419, 
    30.421836419, 30.4211942860001, 30.4204148860001, 30.419268819, 
    30.4138984190001, 30.414127486, 30.4141272190001, 30.4139208190001, 
    30.4136914860001, 30.4132328860001, 30.4131870860001, 30.413255486, 
    30.413599086, 30.4139656190001, 30.4148592190001, 30.4153172860001, 
    30.4157066860001, 30.4160732190001, 30.4168522190001, 30.4181812190001, 
    30.4187540190001, 30.4191664190001, 30.4194868860001, 30.419486686, 
    30.4190734860001, 30.419095886, 30.4192560860001, 30.4195766190001, 
    30.4197596860001, 30.419782019, 30.4199650190001, 30.420125419, 
    30.420720886, 30.420904019, 30.420971219, 30.4211312190001, 
    30.4213832190001, 30.4212222190001, 30.421221819, 30.4214966860001, 
    30.421496486, 30.4213128860001, 30.4205100190001, 30.4200968860001, 
    30.4198442860001, 30.419797886, 30.419660219, 30.4193850190001, 
    30.402990419, 30.404594219, 30.4048692860001, 30.4061982860001, 
    30.4066108860001, 30.407000419, 30.4070920190001, 30.407069086, 
    30.4067478860001, 30.4064038860001, 30.4064726190001, 30.406930819, 
    30.407617686, 30.4083736860001, 30.4086484860001, 30.4092436190001, 
    30.409587286, 30.4103206190001, 30.4106872190001, 30.411832686, 
    30.411970019, 30.395374286, 30.3953510860001, 30.395442686, 
    30.3968164190001, 30.397159619, 30.397938486, 30.398098686, 30.398167019, 
    30.397914219, 30.3976846190001, 30.3971802190001, 30.396996619, 
    30.3968814190001, 30.3963310190001, 30.3956884190001, 30.395023286, 
    30.3944272860001, 30.3934416860001, 30.3917916190001, 30.3915164860001, 
    30.390988819, 30.390713486, 30.3904614190001, 30.3901176190001, 
    30.389522019, 30.388926419, 30.3884908860001, 30.387436419, 
    30.3869550200001, 30.386336086, 30.3860838200001, 30.3860608200001, 
    30.3851434860001, 30.3846158860001, 30.3842950860001, 30.38379102, 
    30.3833326860001, 30.3828512860001, 30.3813154860001, 30.3810176200001, 
    30.3809258200001, 30.378657086, 30.376342886, 30.37519702, 30.373867686, 
    30.373455286, 30.37283662, 30.37201142, 30.3715072200001, 
    30.3854564860001, 30.3852730200001, 30.385043486, 30.3848600200001, 
    30.38456202, 30.38371342, 30.38323202, 30.382613086, 30.381742086, 
    30.380985686, 30.3785562200001, 30.3781206200001, 30.37695102, 
    30.37594202, 30.3751854860001, 30.3743372860001, 30.370623686, 
    30.3691792860001, 30.36842282, 30.3681704860001, 30.3681474860001, 
    30.368559486, 30.369132086, 30.36938422, 30.36968202, 30.3697734200001, 
    30.36952102, 30.369497886, 30.37013862, 30.3706874860001, 30.37116802, 
    30.3708924200001, 30.3709610860001, 30.37242702, 30.372747486, 
    30.3728160200001, 30.3727694200001, 30.3724480860001, 30.3720806200001, 
    30.3715760860001, 30.3715072200001, 30.4119922190001, 30.4120606860001, 
    30.412289619, 30.4128390860001, 30.412976486, 30.412998886, 
    30.4131820860001, 30.4129296190001, 30.4124020190001, 30.412103819, 
    30.4121722190001, 30.4127216860001, 30.4126988190001, 30.411970019, 
    30.411963219, 30.412125486, 30.4121498860001, 30.4119736860001, 
    30.4119922190001, 30.3715072200001, 30.37123222, 30.3706818200001, 
    30.369260486, 30.3689164200001, 30.36834342, 30.36708242, 
    30.3664174200001, 30.3663024200001, 30.3662790860001, 30.366805486, 
    30.36698842, 30.367033486, 30.3669186860001, 30.36641422, 
    30.3659556860001, 30.3651994200001, 30.3644658860001, 30.3641910200001, 
    30.3638474860001, 30.36316062, 30.362702486, 30.362518886, 
    30.3626096200001, 30.362540686, 30.36219642, 30.3619670200001, 
    30.3615772860001, 30.3608438200001, 30.3603622860001, 30.360063886, 
    30.359857086, 30.3598106860001, 30.3599704860001, 30.35987842, 
    30.35836542, 30.3582250200001, 30.3576718200001, 30.35670142, 
    30.35571442, 30.35534102, 30.3543326860001, 30.3534434200001, 
    30.3527990200001, 30.35239482, 30.3522190200001, 30.3519526200001, 
    30.351056086, 30.3469490860001 ;

 flowlines_z = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flowlines_node_count = 25, 4, 20, 23, 7, 4, 62, 5, 9, 48, 41, 44, 44, 21, 
    49, 41, 13, 6, 35, 14 ;

 flowlines_GNIS_NAME =
  "Bull Creek",
  "Bull Creek",
  "Bull Creek",
  "Bull Creek",
  "Bull Creek",
  "Bull Creek",
  "Bull Creek",
  "Bull Creek",
  "Bull Creek",
  "",
  "",
  "",
  "",
  "",
  "West Bull Creek",
  "Cow Fork",
  "",
  "",
  "West Bull Creek",
  "" ;

 catchments_geometry_container = _ ;

 catchments_x = -97.8455203779999, -97.845550745, -97.845238045, 
    -97.8452441169999, -97.844931416, -97.84494963, -97.844636926, 
    -97.8446429969999, -97.8443302909999, -97.844336361, -97.843710948, 
    -97.843717015, -97.8434043079999, -97.843410374, -97.84215954, 
    -97.842171665, -97.841858954, -97.841871077, -97.841558364, 
    -97.841564424, -97.8412517099999, -97.84125777, -97.840319625, 
    -97.840325681, -97.840012965, -97.840025076, -97.839712358, 
    -97.839718412, -97.8394056929999, -97.839411747, -97.839099026, 
    -97.839111131, -97.838798409, -97.8388044609999, -97.838491737, 
    -97.838497788, -97.838185063, -97.8381911129999, -97.837878387, 
    -97.837890484, -97.837577757, -97.837589852, -97.837277122, 
    -97.837283169, -97.836970438, -97.836982529, -97.836669796, 
    -97.836675841, -97.836363107, -97.836369151, -97.83574368, 
    -97.8357557639999, -97.8354430269999, -97.833566602, -97.833572636, 
    -97.8332598979999, -97.833265932, -97.832953192, -97.832959224, 
    -97.832646484, -97.832652515, -97.832339774, -97.8323458039999, 
    -97.8320330609999, -97.832039091, -97.831726347, -97.831732376, 
    -97.831419631, -97.831425659, -97.831112912, -97.831118939, 
    -97.830806192, -97.8308122179999, -97.830186721, -97.830192745, 
    -97.829879996, -97.8298920409999, -97.82957929, -97.8295853119999, 
    -97.8289598059999, -97.8289658259999, -97.8286530729999, -97.828659091, 
    -97.828346337, -97.8283523549999, -97.8277268429999, -97.827732859, 
    -97.8261690739999, -97.826175085, -97.824611293, -97.824617299, 
    -97.82430454, -97.824310544, -97.823997784, -97.824003787, -97.823378264, 
    -97.8233842659999, -97.8230715029999, -97.823077504, -97.822451977, 
    -97.822463974, -97.8227767399999, -97.822782739, -97.822157206, 
    -97.822151208, -97.820900144, -97.8208941509999, -97.820581386, 
    -97.820557416, -97.820244655, -97.820232673, -97.819919914, 
    -97.819913924, -97.819601166, -97.8195951769999, -97.81928242, 
    -97.819276432, -97.818963676, -97.8189576889999, -97.818644934, 
    -97.818603034, -97.818290286, -97.818278317, -97.8179655709999, 
    -97.817959588, -97.817646843, -97.817610949, -97.81729821, 
    -97.8172802669999, -97.816967532, -97.816961552, -97.817274286, 
    -97.817268305, -97.8175810389999, -97.8175750569999, -97.8178877889999, 
    -97.8178818059999, -97.819445462, -97.819439474, -97.8200649349999, 
    -97.820058945, -97.82130986, -97.8213038659999, -97.822867505, 
    -97.822861506, -97.823486959, -97.8234809579999, -97.823793683, 
    -97.8237876809999, -97.824100405, -97.824094402, -97.8244071249999, 
    -97.8244011209999, -97.824713843, -97.8247078379999, -97.8250205589999, 
    -97.825008547, -97.8253212659999, -97.825303245, -97.825615961, 
    -97.8255979369999, -97.82591065, -97.825904641, -97.8265300639999, 
    -97.826524053, -97.827149474, -97.827143461, -97.8274561709999, 
    -97.827450157, -97.8277628659999, -97.8277568509999, -97.828382265, 
    -97.828376248, -97.829001661, -97.8289956419999, -97.8293083469999, 
    -97.8292963069999, -97.82960901, -97.829596968, -97.829909669, 
    -97.829897626, -97.8302103249999, -97.830204302, -97.830517, 
    -97.830510976, -97.8308236729999, -97.830811623, -97.831124318, 
    -97.831112266, -97.8314249589999, -97.831418932, -97.8317316229999, 
    -97.831725596, -97.8320382859999, -97.832032257, -97.832344947, 
    -97.832338917, -97.832651606, -97.832645575, -97.833896324, 
    -97.833890289, -97.834828347, -97.8348223089999, -97.835134994, 
    -97.835128955, -97.8360670069999, -97.8360609649999, -97.836999013, 
    -97.8369929679999, -97.8379310129999, -97.837924965, -97.8382376449999, 
    -97.838550326, -97.8385442759999, -97.838856955, -97.838850904, 
    -97.840101617, -97.840107672, -97.841045709, -97.841051767, 
    -97.841677127, -97.841683188, -97.841995869, -97.84200193, 
    -97.8423146119999, -97.8423206749999, -97.8426333579999, 
    -97.8426394209999, -97.843264789, -97.8432769199999, -97.843589606, 
    -97.843595673, -97.844221047, -97.844227115, -97.844539803, 
    -97.8445519429999, -97.844864633, -97.844876775, -97.845189467, 
    -97.8452016109999, -97.8455143049999, -97.8455203779999, -97.789991152, 
    -97.7899970399999, -97.789684478, -97.7896962519999, -97.789383688, 
    -97.789389574, -97.7890770079999, -97.7890828929999, -97.788770327, 
    -97.788457761, -97.788463644, -97.787838509, -97.78784439, 
    -97.7875318219999, -97.787537702, -97.786599993, -97.78660587, 
    -97.785043016, -97.7850488879999, -97.784736316, -97.7847421869999, 
    -97.784429614, -97.784435484, -97.78412291, -97.7841111719999, 
    -97.784423744, -97.784406135, -97.7847187039999, -97.784712833, 
    -97.785025401, -97.785019529, -97.785332096, -97.785326223, 
    -97.7868890509999, -97.786883173, -97.787508302, -97.787502422, 
    -97.788127549, -97.7881157849999, -97.788428346, -97.788422464, 
    -97.7887350239999, -97.788740908, -97.789991152, -97.775002582, 
    -97.7750084209999, -97.7756336639999, -97.7756395059999, -97.775952128, 
    -97.775957971, -97.776270595, -97.776276439, -97.776589063, 
    -97.7765949079999, -97.7781580339999, -97.778163885, -97.778476511, 
    -97.778482362, -97.7787949889999, -97.778800842, -97.77911347, 
    -97.779119323, -97.779431952, -97.779437807, -97.780375697, 
    -97.780381555, -97.781006817, -97.7810009569999, -97.781938847, 
    -97.7819212589999, -97.782233886, -97.782228022, -97.782540648, 
    -97.782546512, -97.785985404, -97.78599128, -97.786303907, -97.786309784, 
    -97.7869350399999, -97.786940919, -97.787253549, -97.787259429, 
    -97.787572059, -97.7875779399999, -97.787890572, -97.787896454, 
    -97.7882090859999, -97.788214969, -97.788527603, -97.7885334869999, 
    -97.7919724609999, -97.7919665649999, -97.792279198, -97.792273301, 
    -97.7925859329999, -97.792580035, -97.792892665, -97.792886767, 
    -97.793199396, -97.793193496, -97.794131382, -97.7941254789999, 
    -97.795688615, -97.795694523, -97.796319779, -97.796325689, 
    -97.796638318, -97.7966324069999, -97.796945035, -97.797257663, 
    -97.797263576, -97.7985140919999, -97.798826721, -97.7988503939999, 
    -97.798537761, -97.798596937, -97.798284294, -97.798307961, 
    -97.798620608, -97.798662035, -97.798974689, -97.798992447, 
    -97.799305105, -97.7993465489999, -97.799033884, -97.7990457229999, 
    -97.7987330559999, -97.798738975, -97.7984263069999, -97.7984322249999, 
    -97.798119556, -97.798125473, -97.7984381429999, -97.79844406, 
    -97.799069402, -97.7990812419999, -97.799706588, -97.7997125099999, 
    -97.800025184, -97.8000311069999, -97.800343782, -97.800349706, 
    -97.8009750579999, -97.800980984, -97.801293661, -97.801305516, 
    -97.8016181949999, -97.801624123, -97.801936803, -97.801942732, 
    -97.802255413, -97.802261344, -97.8025740259999, -97.802579957, 
    -97.80289264, -97.802910438, -97.8032231239999, -97.8032349919999, 
    -97.802922304, -97.802946036, -97.802633344, -97.802639276, 
    -97.802326583, -97.8023325139999, -97.802019819, -97.8020257489999, 
    -97.8017130539999, -97.8017189829999, -97.801406287, -97.801412215, 
    -97.801099517, -97.801105445, -97.800792746, -97.800798672, 
    -97.7989224739999, -97.798916554, -97.797978458, -97.797972541, 
    -97.7973471449999, -97.797341231, -97.797028534, -97.79702262, 
    -97.796397228, -97.796391317, -97.794827841, -97.794821935, 
    -97.793883853, -97.7938897559999, -97.793264365, -97.793270267, 
    -97.792332177, -97.792326279, -97.792013584, -97.792007687, 
    -97.791694992, -97.791689096, -97.791063709, -97.791057815, -97.79043243, 
    -97.790426538, -97.789801155, -97.789795265, -97.789482575, 
    -97.789470797, -97.789158109, -97.789134559, -97.788821874, 
    -97.788786556, -97.788473878, -97.788467993, -97.787842638, 
    -97.7878367549999, -97.787524078, -97.7875181969999, -97.787205521, 
    -97.78719964, -97.786574291, -97.786568412, -97.785630392, 
    -97.7856186399999, -97.785305969, -97.785300094, -97.784674753, 
    -97.78466888, -97.784356211, -97.784350339, -97.783725002, -97.783719133, 
    -97.78121779, -97.7812119289999, -97.780899262, -97.7808934019999, 
    -97.778079406, -97.775890741, -97.775884897, -97.775259566, 
    -97.775253725, -97.7749410599999, -97.77493522, -97.774309893, 
    -97.774304054, -97.773991392, -97.773985554, -97.773672893, 
    -97.773667057, -97.7733543959999, -97.773348561, -97.773035901, 
    -97.773030067, -97.771779432, -97.7717736019999, -97.771148286, 
    -97.771142459, -97.770517145, -97.770505494, -97.7701928389999, 
    -97.770187014, -97.76987436, -97.769862713, -97.769550061, -97.769538417, 
    -97.769225767, -97.769219946, -97.7689072969999, -97.768901477, 
    -97.769214124, -97.769208303, -97.7698335969999, -97.769821951, 
    -97.7701345949999, -97.770128771, -97.7704414149999, -97.7704239399999, 
    -97.7707365799999, -97.770719102, -97.77103174, -97.771020086, 
    -97.771332721, -97.771315237, -97.77162787, -97.7716103829999, 
    -97.7719230119999, -97.771917183, -97.772229811, -97.77222398, 
    -97.772536607, -97.772530775, -97.772843401, -97.7728375679999, 
    -97.773150193, -97.773144359, -97.773456983, -97.773451148, 
    -97.774076394, -97.774070557, -97.7746958, -97.774689961, -97.775002582, 
    -97.788770327, -97.788782095, -97.789407232, -97.789413118, 
    -97.789725687, -97.789731574, -97.790044145, -97.7900500329999, 
    -97.7903626039999, -97.790368493, -97.790993638, -97.790999529, 
    -97.7913121019999, -97.791335673, -97.79164825, -97.7916777189999, 
    -97.7919903009999, -97.792002091, -97.7923146749999, -97.7923264679999, 
    -97.7926390539999, -97.7926862319999, -97.792998827, -97.7930047249999, 
    -97.793317321, -97.79332322, -97.7936358169999, -97.793647618, 
    -97.793960216, -97.793977922, -97.794290523, -97.794320038, 
    -97.794632645, -97.794644453, -97.794957061, -97.794986588, 
    -97.795299202, -97.795311014, -97.79562363, -97.795635445, -97.795948063, 
    -97.7959598799999, -97.7962725, -97.79627841, -97.796903652, 
    -97.796945035, -97.7966324069999, -97.796638318, -97.796325689, 
    -97.796319779, -97.795694523, -97.795688615, -97.7941254789999, 
    -97.794131382, -97.793193496, -97.793199396, -97.792886767, 
    -97.792892665, -97.792580035, -97.7925859329999, -97.792273301, 
    -97.792279198, -97.7919665649999, -97.7919724609999, -97.7885334869999, 
    -97.788527603, -97.788214969, -97.7882090859999, -97.787896454, 
    -97.787890572, -97.7875779399999, -97.787572059, -97.787259429, 
    -97.787253549, -97.786940919, -97.7869350399999, -97.786309784, 
    -97.786303907, -97.78599128, -97.785985404, -97.782546512, -97.782540648, 
    -97.782228022, -97.782233886, -97.7819212589999, -97.781938847, 
    -97.7810009569999, -97.781006817, -97.780381555, -97.780375697, 
    -97.779437807, -97.779431952, -97.779119323, -97.77911347, -97.778800842, 
    -97.7787949889999, -97.778482362, -97.778476511, -97.778163885, 
    -97.7781580339999, -97.7765949079999, -97.776589063, -97.776276439, 
    -97.776270595, -97.775957971, -97.775952128, -97.7756395059999, 
    -97.7756336639999, -97.7750084209999, -97.775002582, -97.774985063, 
    -97.774672445, -97.774643253, -97.774955865, -97.7749208289999, 
    -97.775233436, -97.775215915, -97.775210075, -97.775522677, 
    -97.775516836, -97.775829437, -97.775817753, -97.7761303509999, 
    -97.776118665, -97.776431262, -97.776419574, -97.776732169, 
    -97.776726324, -97.777976697, -97.7779708479999, -97.778908625, 
    -97.7789144769999, -97.779539663, -97.779545517, -97.780170706, 
    -97.780176562, -97.780489157, -97.7804833, -97.7807958939999, 
    -97.780778319, -97.78109091, -97.781067473, -97.7813800599999, 
    -97.7813742, -97.781686786, -97.781680925, -97.781993509, -97.781981785, 
    -97.782294368, -97.782282642, -97.7825952219999, -97.7825893579999, 
    -97.782901938, -97.782896073, -97.7832086509999, -97.783202785, 
    -97.7835153619999, -97.783509495, -97.783822072, -97.7838162039999, 
    -97.784128779, -97.78412291, -97.784435484, -97.784429614, 
    -97.7847421869999, -97.784736316, -97.7850488879999, -97.785043016, 
    -97.78660587, -97.786599993, -97.787537702, -97.7875318219999, 
    -97.78784439, -97.787838509, -97.788463644, -97.788457761, -97.788770327, 
    -97.7701928389999, -97.769880184, -97.76987436, -97.770187014, 
    -97.7701928389999, -97.7701928389999, -97.770505494, -97.770517145, 
    -97.771142459, -97.771148286, -97.7717736019999, -97.771779432, 
    -97.773030067, -97.773035901, -97.773348561, -97.7733543959999, 
    -97.773667057, -97.773672893, -97.773985554, -97.773991392, 
    -97.774304054, -97.774309893, -97.77493522, -97.7749410599999, 
    -97.775253725, -97.775259566, -97.775884897, -97.775890741, 
    -97.778079406, -97.778085257, -97.775896584, -97.7759024279999, 
    -97.775589759, -97.775595602, -97.775282932, -97.775306299, 
    -97.774993625, -97.7749994659999, -97.774686791, -97.7746926299999, 
    -97.774379954, -97.774385793, -97.774073116, -97.7740789539999, 
    -97.773766275, -97.773807133, -97.773494448, -97.773500284, -97.77350612, 
    -97.772880745, -97.772886579, -97.77257389, -97.772579723, 
    -97.7719543439999, -97.7719601749999, -97.771647484, -97.771653314, 
    -97.771340622, -97.7713464509999, -97.770408372, -97.770414198, 
    -97.76978881, -97.769777163, -97.7694644699999, -97.769423712, 
    -97.769111027, -97.769105205, -97.768792521, -97.768786701, 
    -97.7684740179999, -97.7684565599999, -97.76876924, -97.7687168589999, 
    -97.769029529, -97.769017887, -97.7693305559999, -97.769301446, 
    -97.76961411, -97.769596642, -97.769909302, -97.769886007, -97.770198663, 
    -97.7701928389999, -97.809080509, -97.809086464, -97.808773684, 
    -97.808779638, -97.808466857, -97.808490669, -97.808177884, 
    -97.8081897879999, -97.807877001, -97.807906757, -97.807593964, 
    -97.807599915, -97.8072871209999, -97.8072930709999, -97.806667481, 
    -97.8066734289999, -97.8063606329999, -97.806366579, -97.806053783, 
    -97.806059728, -97.8057469299999, -97.805752874, -97.805440076, 
    -97.805422246, -97.805735042, -97.805717209, -97.8060300019999, 
    -97.8060240569999, -97.8063368479999, -97.8063130639999, -97.806625852, 
    -97.806608011, -97.8069207949999, -97.806897004, -97.807209784, 
    -97.807203836, -97.809080509, -97.778079406, -97.7808934019999, 
    -97.780899262, -97.7812119289999, -97.78121779, -97.783719133, 
    -97.783725002, -97.784350339, -97.784356211, -97.78466888, -97.784674753, 
    -97.785300094, -97.785305969, -97.7856186399999, -97.785630392, 
    -97.786568412, -97.786574291, -97.78719964, -97.787205521, 
    -97.7875181969999, -97.787524078, -97.7878367549999, -97.787842638, 
    -97.788467993, -97.788473878, -97.788786556, -97.788821874, 
    -97.789134559, -97.789158109, -97.789470797, -97.789482575, 
    -97.789795265, -97.789801155, -97.790426538, -97.79043243, -97.791057815, 
    -97.791063709, -97.791689096, -97.791694992, -97.792007687, 
    -97.792013584, -97.792326279, -97.792332177, -97.793270267, 
    -97.793264365, -97.7938897559999, -97.793883853, -97.794821935, 
    -97.794827841, -97.796391317, -97.796397228, -97.79702262, -97.797028534, 
    -97.797341231, -97.7973471449999, -97.797972541, -97.797978458, 
    -97.798916554, -97.7989224739999, -97.800798672, -97.800804598, 
    -97.8011172989999, -97.801129153, -97.8014418559999, -97.801453712, 
    -97.801766417, -97.8017782759999, -97.802403689, -97.802409621, 
    -97.803035036, -97.8030409689999, -97.803979095, -97.803985031, 
    -97.80492316, -97.804929099, -97.80524181, -97.805247751, -97.805560462, 
    -97.805566404, -97.805879116, -97.805885059, -97.806510486, 
    -97.806516431, -97.8068291449999, -97.806835092, -97.807460522, 
    -97.8074664709999, -97.8077791869999, -97.807785136, -97.8080978529999, 
    -97.808103804, -97.808416522, -97.8084224739999, -97.808735193, 
    -97.8087411449999, -97.809366586, -97.80937254, -97.809685261, 
    -97.809691217, -97.810003939, -97.8100098959999, -97.810322619, 
    -97.810334535, -97.8106472599999, -97.810653219, -97.810965945, 
    -97.810971905, -97.811284632, -97.811290594, -97.8116033219999, 
    -97.811609284, -97.811922013, -97.8119279759999, -97.812240706, 
    -97.812246671, -97.8131848639999, -97.813190831, -97.813503563, 
    -97.8135154999999, -97.8141409679999, -97.814146939, -97.815710613, 
    -97.815716589, -97.816967532, -97.8172802669999, -97.81729821, 
    -97.817610949, -97.817646843, -97.817959588, -97.8179655709999, 
    -97.818278317, -97.818290286, -97.818603034, -97.818644934, 
    -97.818332179, -97.818344149, -97.8177186349999, -97.8177306009999, 
    -97.817417841, -97.817435788, -97.8171230249999, -97.817129006, 
    -97.815565189, -97.8155711649999, -97.814945635, -97.814951609, 
    -97.8146388439999, -97.814644817, -97.813706516, -97.813712486, 
    -97.813399718, -97.813411656, -97.812786116, -97.812792083, 
    -97.811853769, -97.811865697, -97.811552923, -97.811564849, 
    -97.8106265229999, -97.8106324829999, -97.810319706, -97.809694153, 
    -97.8097001099999, -97.809387332, -97.809393288, -97.809080509, 
    -97.807203836, -97.807209784, -97.806897004, -97.8069207949999, 
    -97.806608011, -97.806625852, -97.8063130639999, -97.8063368479999, 
    -97.8060240569999, -97.8060300019999, -97.805717209, -97.805735042, 
    -97.805422246, -97.805440076, -97.805446019, -97.805133219, 
    -97.8051391609999, -97.8048263599999, -97.8048382429999, -97.80452544, 
    -97.804543261, -97.8048560669999, -97.804873892, -97.805186701, 
    -97.805216415, -97.8055292289999, -97.805558949, -97.805246129, 
    -97.805275845, -97.8049630199999, -97.804980847, -97.805293675, 
    -97.805311505, -97.8056243359999, -97.805660003, -97.80597284, 
    -97.806014461, -97.805701617, -97.805713507, -97.805400661, 
    -97.8054244369999, -97.8051115869999, -97.805129417, -97.80544227, 
    -97.805460103, -97.80577296, -97.8057848509999, -97.806097709, 
    -97.806115549, -97.806428411, -97.8064819419999, -97.806794813, 
    -97.806806711, -97.807119584, -97.807155286, -97.807468165, 
    -97.807486019, -97.807798901, -97.807810806, -97.8081236899999, 
    -97.808129644, -97.808442529, -97.8084484839999, -97.80876137, 
    -97.808767326, -97.809080213, -97.8090861699999, -97.8093990579999, 
    -97.809405016, -97.809717905, -97.809723864, -97.810349644, 
    -97.810361566, -97.8106744579999, -97.810680421, -97.810993313, 
    -97.810999277, -97.8113121709999, -97.811318135, -97.8116310299999, 
    -97.8116369959999, -97.811949892, -97.811955858, -97.8125816519999, 
    -97.812587621, -97.809771538, -97.809777498, -97.809151699, 
    -97.8091457419999, -97.808207046, -97.808213001, -97.8069614029999, 
    -97.8069673529999, -97.8063415509999, -97.806335603, -97.8057098039999, 
    -97.80571575, -97.803838344, -97.803844284, -97.801653969, -97.801648036, 
    -97.801022234, -97.801016303, -97.7991388999999, -97.799132976, 
    -97.797255578, -97.797261496, -97.79538409, -97.795378178, -97.794439478, 
    -97.794433569, -97.793807771, -97.793801864, -97.792863169, 
    -97.792857265, -97.7925443679999, -97.792538465, -97.791912673, 
    -97.7919067719999, -97.791593877, -97.7915879769999, -97.790962189, 
    -97.790956291, -97.790643398, -97.790637502, -97.790324609, 
    -97.790318714, -97.789692931, -97.789687038, -97.789374148, 
    -97.789368256, -97.788742477, -97.788736587, -97.788423698, 
    -97.788417809, -97.7881049219999, -97.788081371, -97.7877684869999, 
    -97.787744941, -97.7874320609999, -97.787420291, -97.7871074129999, 
    -97.787101529, -97.786788653, -97.786776886, -97.786464012, 
    -97.786458129, -97.7861452559999, -97.786133494, -97.785820623, 
    -97.7858147429999, -97.7855018719999, -97.785490114, -97.785177246, 
    -97.785171368, -97.784858501, -97.7848526239999, -97.7845397579999, 
    -97.7845338819999, -97.7842210169999, -97.7842151419999, 
    -97.7832765489999, -97.783270678, -97.782957814, -97.782963685, 
    -97.782337956, -97.782332087, -97.782019224, -97.782025091, 
    -97.7813993619999, -97.7814052269999, -97.781092362, -97.781098226, 
    -97.7804724919999, -97.780478355, -97.780165487, -97.780171348, 
    -97.77954561, -97.7795514699999, -97.778612859, -97.778607003, 
    -97.778294134, -97.778288279, -97.777662542, -97.777656689, 
    -97.777343822, -97.77733797, -97.777025104, -97.776712238, -97.776706388, 
    -97.776393522, -97.776387673, -97.776074809, -97.776068961, 
    -97.775443235, -97.775437389, -97.774811664, -97.774805821, 
    -97.774492959, -97.774487117, -97.773861396, -97.7738555559999, 
    -97.7735426959999, -97.773536857, -97.77291114, -97.772905303, 
    -97.7722795879999, -97.772273753, -97.7719608959999, -97.771955062, 
    -97.771329351, -97.771323519, -97.7706978099999, -97.77069198, 
    -97.770379126, -97.770373297, -97.769747592, -97.769741765, 
    -97.769116062, -97.769110237, -97.768797386, -97.768791563, 
    -97.768165863, -97.768160042, -97.767534344, -97.767528525, 
    -97.767215677, -97.767209859, -97.766584165, -97.766578349, 
    -97.766566717, -97.7668795599999, -97.766867926, -97.7671807679999, 
    -97.76717495, -97.76748779, -97.7674819709999, -97.767794811, 
    -97.767788991, -97.768101829, -97.768090187, -97.768403024, 
    -97.768397202, -97.7687100369999, -97.768704214, -97.769017048, 
    -97.7690112239999, -97.7693240579999, -97.769312408, -97.7696252389999, 
    -97.769607761, -97.769920589, -97.769914762, -97.7702275889999, 
    -97.770221761, -97.770534587, -97.77052293, -97.770835753, 
    -97.7708299239999, -97.771142746, -97.771136916, -97.771449737, 
    -97.771443905, -97.771756726, -97.771750893, -97.772063713, 
    -97.772057879, -97.772370697, -97.772364863, -97.773303314, 
    -97.773297477, -97.773610293, -97.773604454, -97.773917269, 
    -97.773911429, -97.7761011269999, -97.7760952799999, -97.777972156, 
    -97.777966303, -97.778279115, -97.778273261, -97.778898881, 
    -97.778887169, -97.779199978, -97.779182407, -97.779495212, 
    -97.779465922, -97.7797787219999, -97.7797611459999, -97.780073943, 
    -97.7800622239999, -97.779749429, -97.779725995, -97.780038786, 
    -97.780027067, -97.780339855, -97.780322274, -97.780009489, 
    -97.780003629, -97.7796908449999, -97.7796849869999, -97.779372203, 
    -97.779366346, -97.779679129, -97.779667412, -97.779980193, 
    -97.779927462, -97.7796146909999, -97.779608834, -97.7792960639999, 
    -97.779290207, -97.778977438, -97.7789715819999, -97.778658814, 
    -97.7786471049999, -97.778334339, -97.778328486, -97.7777029549999, 
    -97.777697104, -97.77738434, -97.77737849, -97.777065726, -97.777048179, 
    -97.7773609389999, -97.777325839, -97.777013085, -97.777001388, 
    -97.776688636, -97.7766710929999, -97.776358344, -97.776317419, 
    -97.7760046769999, -97.7759520709999, -97.7762648039999, -97.776229729, 
    -97.775917002, -97.775887779, -97.775575058, -97.775557528, 
    -97.7752448099999, -97.775203914, -97.774891203, -97.774826954, 
    -97.775139654, -97.775127971, -97.775440668, -97.775423141, 
    -97.775735835, -97.775706618, -97.775393929, -97.775388086, 
    -97.775075398, -97.7750695569999, -97.7738188069999, -97.7738129699999, 
    -97.773500284, -97.773494448, -97.773807133, -97.773766275, 
    -97.7740789539999, -97.774073116, -97.774385793, -97.774379954, 
    -97.7746926299999, -97.774686791, -97.7749994659999, -97.774993625, 
    -97.775306299, -97.775282932, -97.775595602, -97.775589759, 
    -97.7759024279999, -97.775896584, -97.778085257, -97.778079406, 
    -97.810319706, -97.810373338, -97.810686124, -97.810721886, 
    -97.810409094, -97.8104210129999, -97.810432933, -97.810120136, 
    -97.810126095, -97.8098132979999, -97.80980734, -97.809494544, 
    -97.809488587, -97.809175792, -97.809169837, -97.808544248, 
    -97.8085382949999, -97.8079127079999, -97.807906757, -97.807877001, 
    -97.8081897879999, -97.808177884, -97.808490669, -97.808466857, 
    -97.808779638, -97.808773684, -97.809086464, -97.809080509, 
    -97.809393288, -97.809387332, -97.8097001099999, -97.809694153, 
    -97.810319706, -97.818644934, -97.8189576889999, -97.818963676, 
    -97.819276432, -97.81928242, -97.8195951769999, -97.819601166, 
    -97.819913924, -97.819919914, -97.820232673, -97.820244655, 
    -97.820557416, -97.820581386, -97.8208941509999, -97.820900144, 
    -97.822151208, -97.822157206, -97.822782739, -97.822788739, 
    -97.823101507, -97.823107508, -97.823420277, -97.823426279, 
    -97.8237390479999, -97.8237450509999, -97.824057822, -97.824063826, 
    -97.824376598, -97.8243826029999, -97.824695376, -97.8247013819999, 
    -97.825014156, -97.825020163, -97.825332938, -97.825356971, -97.82566975, 
    -97.825681769, -97.825687779, -97.825374997, -97.8253810049999, 
    -97.825068222, -97.82507423, -97.824761446, -97.8247674529999, 
    -97.824454668, -97.824460673, -97.823835101, -97.8238411039999, 
    -97.8219643799999, -97.8219703779999, -97.821344801, -97.821350796, 
    -97.820725217, -97.82073121, -97.820105629, -97.82011162, -97.818860452, 
    -97.81886644, -97.8169896809999, -97.8169837, -97.81323019, 
    -97.813224221, -97.8129114289999, -97.812917397, -97.810727847, 
    -97.810733807, -97.8104210129999, -97.810409094, -97.810721886, 
    -97.810686124, -97.810373338, -97.810319706, -97.8106324829999, 
    -97.8106265229999, -97.811564849, -97.811552923, -97.811865697, 
    -97.811853769, -97.812792083, -97.812786116, -97.813411656, 
    -97.813399718, -97.813712486, -97.813706516, -97.814644817, 
    -97.8146388439999, -97.814951609, -97.814945635, -97.8155711649999, 
    -97.815565189, -97.817129006, -97.8171230249999, -97.817435788, 
    -97.817417841, -97.8177306009999, -97.8177186349999, -97.818344149, 
    -97.818332179, -97.818644934, -97.7685872439999, -97.768899837, 
    -97.768905656, -97.769530843, -97.769536664, -97.770474447, 
    -97.7704802709999, -97.770792866, -97.770798692, -97.771111288, 
    -97.771122941, -97.771435539, -97.771441367, -97.772379164, 
    -97.772384995, -97.772697595, -97.772703427, -97.773328629, 
    -97.773334463, -97.7742722689999, -97.7742781059999, -97.775215915, 
    -97.775233436, -97.7749208289999, -97.774955865, -97.774643253, 
    -97.774672445, -97.774985063, -97.775002582, -97.774689961, -97.7746958, 
    -97.774070557, -97.774076394, -97.773451148, -97.773456983, 
    -97.773144359, -97.773150193, -97.7728375679999, -97.772843401, 
    -97.772530775, -97.772536607, -97.77222398, -97.772229811, -97.771917183, 
    -97.7719230119999, -97.7716103829999, -97.77162787, -97.771315237, 
    -97.771332721, -97.771020086, -97.77103174, -97.770719102, 
    -97.7707365799999, -97.7704239399999, -97.7704414149999, -97.770128771, 
    -97.7701345949999, -97.769821951, -97.7698335969999, -97.769208303, 
    -97.769214124, -97.768901477, -97.7689072969999, -97.769219946, 
    -97.769225767, -97.769538417, -97.769550061, -97.769862713, -97.76987436, 
    -97.769880184, -97.7701928389999, -97.770198663, -97.769886007, 
    -97.769909302, -97.769596642, -97.76961411, -97.769301446, 
    -97.7693305559999, -97.769017887, -97.769029529, -97.7687168589999, 
    -97.76876924, -97.7684565599999, -97.7684740179999, -97.768786701, 
    -97.768792521, -97.769105205, -97.769111027, -97.769423712, 
    -97.7694644699999, -97.769777163, -97.76978881, -97.769476116, 
    -97.7694819389999, -97.769169244, -97.7691750659999, -97.76886237, 
    -97.76886819, -97.768555493, -97.768561313, -97.7682486149999, 
    -97.7682777099999, -97.7679650059999, -97.7679766429999, -97.767663937, 
    -97.7676697539999, -97.767044341, -97.767050156, -97.766737448, 
    -97.7667723329999, -97.767085047, -97.76711994, -97.76680722, 
    -97.7668188499999, -97.766506127, -97.766529382, -97.766842109, 
    -97.766859553, -97.767172283, -97.767183915, -97.767496646, 
    -97.767514098, -97.767826832, -97.7678442869999, -97.7681570239999, 
    -97.7682152199999, -97.7685279679999, -97.76854543, -97.7682326789999, 
    -97.768244319, -97.767931566, -97.767937385, -97.767624631, 
    -97.767630449, -97.767317694, -97.767323511, -97.7670107549999, 
    -97.7670340189999, -97.767346779, -97.767364231, -97.7676769939999, 
    -97.767694449, -97.768007215, -97.768018854, -97.7683316229999, 
    -97.768354905, -97.768667678, -97.768679321, -97.768992096, 
    -97.7690037409999, -97.769316518, -97.769328166, -97.769015387, 
    -97.769032856, -97.7693456379999, -97.7693572859999, -97.76967007, 
    -97.7696875459999, -97.7700003319999, -97.7700119849999, -97.769699196, 
    -97.769734149, -97.7700469439999, -97.7700527709999, -97.7703655669999, 
    -97.770371395, -97.770684192, -97.770690021, -97.771002819, 
    -97.771014478, -97.7713272779999, -97.771344771, -97.771657574, 
    -97.7716809029999, -97.7719937099999, -97.771999544, -97.772312352, 
    -97.772318186, -97.772630995, -97.7726368309999, -97.772949641, 
    -97.772955477, -97.7732682879999, -97.773274126, -97.7735869379999, 
    -97.773592777, -97.77390559, -97.773911429, -97.773917269, -97.773604454, 
    -97.773610293, -97.773297477, -97.773303314, -97.772364863, 
    -97.772370697, -97.772057879, -97.772063713, -97.771750893, 
    -97.771756726, -97.771443905, -97.771449737, -97.771136916, 
    -97.771142746, -97.7708299239999, -97.770835753, -97.77052293, 
    -97.770534587, -97.770221761, -97.7702275889999, -97.769914762, 
    -97.769920589, -97.769607761, -97.7696252389999, -97.769312408, 
    -97.7693240579999, -97.7690112239999, -97.769017048, -97.768704214, 
    -97.7687100369999, -97.768397202, -97.768403024, -97.768090187, 
    -97.768101829, -97.767788991, -97.767794811, -97.7674819709999, 
    -97.76748779, -97.76717495, -97.7671807679999, -97.766867926, 
    -97.7668795599999, -97.766566717, -97.766578349, -97.765952657, 
    -97.7659468429999, -97.7656339979999, -97.765628185, -97.765002497, 
    -97.764996686, -97.764371, -97.764365191, -97.7640523489999, 
    -97.764046541, -97.763420859, -97.763415054, -97.762789373, -97.76278357, 
    -97.762470731, -97.762464928, -97.761839252, -97.761833451, 
    -97.761207777, -97.761201978, -97.760576306, -97.76057051, -97.759944839, 
    -97.759939045, -97.759626211, -97.7596204179999, -97.758994751, 
    -97.75898896, -97.758363295, -97.758357506, -97.758044675, 
    -97.7580388869999, -97.757413226, -97.75740744, -97.756781781, 
    -97.756775998, -97.756463169, -97.756457386, -97.7558317309999, 
    -97.755825951, -97.755200298, -97.755194519, -97.7548816939999, 
    -97.7548759159999, -97.754250267, -97.7542444919999, -97.753618844, 
    -97.753613071, -97.7529874259999, -97.752981655, -97.752668833, 
    -97.7526630629999, -97.752037421, -97.752031654, -97.7514060139999, 
    -97.751400248, -97.7510874289999, -97.751081665, -97.750768847, 
    -97.750763083, -97.750137449, -97.750131688, -97.749506056, 
    -97.749500296, -97.749187481, -97.7491817229999, -97.748556095, 
    -97.748544582, -97.74823177, -97.74822026, -97.74790745, -97.747901696, 
    -97.7475888869999, -97.747577381, -97.747264574, -97.747253071, 
    -97.746940266, -97.746905762, -97.746592963, -97.746552717, 
    -97.746239926, -97.746205437, -97.745892651, -97.7458696639999, 
    -97.7455568829999, -97.745539645, -97.745226867, -97.745203889, 
    -97.745516663, -97.745510918, -97.745198144, -97.745163678, 
    -97.744850911, -97.744839425, -97.74452666, -97.744486466, -97.744799224, 
    -97.7447762529999, -97.745089007, -97.745071776, -97.745384526, 
    -97.745378782, -97.745066032, -97.745060289, -97.745373037, 
    -97.745350059, -97.7456628039999, -97.7456455669999, -97.7459583089999, 
    -97.745946816, -97.7462595549999, -97.746248061, -97.746560798, 
    -97.746549301, -97.746862036, -97.746850538, -97.747163271, 
    -97.7471517709999, -97.747464502, -97.747452999, -97.747765728, 
    -97.7477599759999, -97.748072704, -97.748061198, -97.748373923, 
    -97.748362415, -97.7486751389999, -97.748669384, -97.748982106, 
    -97.74897635, -97.749289072, -97.749283315, -97.749596035, 
    -97.7495499729999, -97.74923726, -97.749225747, -97.748913037, 
    -97.7489015259999, -97.748588818, -97.7485830639999, -97.748270357, 
    -97.74825885, -97.747946145, -97.747940393, -97.747627689, -97.747621938, 
    -97.747309235, -97.747303485, -97.7469907829999, -97.746979285, 
    -97.746666585, -97.746660837, -97.746348138, -97.746342391, 
    -97.746029693, -97.746023947, -97.7457112499999, -97.745699761, 
    -97.745387066, -97.745381322, -97.745068628, -97.7450571429999, 
    -97.745369835, -97.745364092, -97.745676783, -97.745665294, 
    -97.7459779819999, -97.745955001, -97.745642316, -97.7456308279999, 
    -97.7453181449999, -97.745300916, -97.745613595, -97.745602107, 
    -97.745914785, -97.74590904, -97.746221716, -97.746210224, -97.746522898, 
    -97.746505658, -97.746818329, -97.74678959, -97.7471022559999, 
    -97.74708501, -97.747397673, -97.747391923, -97.747704585, 
    -97.7476988339999, -97.748011495, -97.748005743, -97.748318403, 
    -97.748312651, -97.748625309, -97.7486195559999, -97.748932213, 
    -97.7489207039999, -97.7492333599999, -97.7492276039999, -97.749540258, 
    -97.749534502, -97.7498471549999, -97.74983564, -97.750148291, 
    -97.750142533, -97.750455183, -97.750449424, -97.750762073, 
    -97.750756312, -97.7510689599999, -97.751063199, -97.751375846, 
    -97.751370084, -97.751682729, -97.751676966, -97.7526149, -97.752609134, 
    -97.753547065, -97.753541295, -97.754479223, -97.754473451, 
    -97.754786092, -97.754780318, -97.755092959, -97.7550814099999, 
    -97.755394048, -97.7553882719999, -97.75570091, -97.7556893569999, 
    -97.7560019919999, -97.7559962139999, -97.7563088479999, 
    -97.7562972919999, -97.756609924, -97.7566041439999, -97.756916775, 
    -97.756905214, -97.757217843, -97.757212062, -97.75752469, -97.757518907, 
    -97.757831534, -97.757825751, -97.758763627, -97.758757841, -97.75938309, 
    -97.759377301, -97.759689925, -97.759684135, -97.76030938, 
    -97.7603035879999, -97.76061621, -97.760610417, -97.7609230369999, 
    -97.760917244, -97.761229863, -97.761206686, -97.7608940709999, 
    -97.7608708989999, -97.761183509, -97.761171921, -97.76148453, 
    -97.76147294, -97.761785547, -97.7617797509999, -97.7624049619999, 
    -97.762399164, -97.762711768, -97.762705969, -97.763018573, 
    -97.763012773, -97.763637977, -97.7636321749999, -97.7648825799999, 
    -97.764876774, -97.7670649729999, -97.76705916, -97.767371759, 
    -97.7673659449999, -97.767678543, -97.767672727, -97.7679853239999, 
    -97.7679795079999, -97.768292103, -97.7682746519999, -97.7685872439999, 
    -97.773500284, -97.7738129699999, -97.7738188069999, -97.7750695569999, 
    -97.775075398, -97.775388086, -97.775393929, -97.775706618, 
    -97.775735835, -97.775423141, -97.775440668, -97.775127971, 
    -97.775139654, -97.774826954, -97.774891203, -97.775203914, 
    -97.7752448099999, -97.775557528, -97.775575058, -97.775887779, 
    -97.775917002, -97.776229729, -97.7762648039999, -97.7759520709999, 
    -97.7760046769999, -97.776317419, -97.776358344, -97.7766710929999, 
    -97.776688636, -97.777001388, -97.777013085, -97.777325839, 
    -97.7773609389999, -97.777048179, -97.777065726, -97.77737849, 
    -97.77738434, -97.777697104, -97.7777029549999, -97.778328486, 
    -97.778334339, -97.7786471049999, -97.778658814, -97.7789715819999, 
    -97.778977438, -97.779290207, -97.7792960639999, -97.779608834, 
    -97.7796146909999, -97.779927462, -97.779980193, -97.779667412, 
    -97.779679129, -97.779366346, -97.779372203, -97.7796849869999, 
    -97.7796908449999, -97.780003629, -97.780009489, -97.780322274, 
    -97.780339855, -97.780027067, -97.780038786, -97.779725995, 
    -97.779749429, -97.7800622239999, -97.780073943, -97.7797611459999, 
    -97.7797787219999, -97.779465922, -97.779495212, -97.779182407, 
    -97.779199978, -97.778887169, -97.778898881, -97.778273261, 
    -97.778279115, -97.777966303, -97.777972156, -97.7760952799999, 
    -97.7761011269999, -97.773911429, -97.77390559, -97.773592777, 
    -97.7735869379999, -97.773274126, -97.7732682879999, -97.772955477, 
    -97.772949641, -97.7726368309999, -97.772630995, -97.772318186, 
    -97.772312352, -97.771999544, -97.7719937099999, -97.7716809029999, 
    -97.771657574, -97.771344771, -97.7713272779999, -97.771014478, 
    -97.771002819, -97.770690021, -97.770684192, -97.770371395, 
    -97.7703655669999, -97.7700527709999, -97.7700469439999, -97.769734149, 
    -97.769699196, -97.7700119849999, -97.7700003319999, -97.7696875459999, 
    -97.76967007, -97.7693572859999, -97.7693456379999, -97.769032856, 
    -97.769015387, -97.769328166, -97.769316518, -97.7690037409999, 
    -97.768992096, -97.768679321, -97.768667678, -97.768354905, 
    -97.7683316229999, -97.768018854, -97.768007215, -97.767694449, 
    -97.7676769939999, -97.767364231, -97.767346779, -97.7670340189999, 
    -97.7670107549999, -97.767323511, -97.767317694, -97.767630449, 
    -97.767624631, -97.767937385, -97.767931566, -97.768244319, 
    -97.7682326789999, -97.76854543, -97.7685279679999, -97.7682152199999, 
    -97.7681570239999, -97.7678442869999, -97.767826832, -97.767514098, 
    -97.767496646, -97.767183915, -97.767172283, -97.766859553, 
    -97.766842109, -97.766529382, -97.766506127, -97.7668188499999, 
    -97.76680722, -97.76711994, -97.767085047, -97.7667723329999, 
    -97.766737448, -97.767050156, -97.767044341, -97.7676697539999, 
    -97.767663937, -97.7679766429999, -97.7679650059999, -97.7682777099999, 
    -97.7682486149999, -97.768561313, -97.768555493, -97.76886819, 
    -97.76886237, -97.7691750659999, -97.769169244, -97.7694819389999, 
    -97.769476116, -97.76978881, -97.770414198, -97.770408372, 
    -97.7713464509999, -97.771340622, -97.771653314, -97.771647484, 
    -97.7719601749999, -97.7719543439999, -97.772579723, -97.77257389, 
    -97.772886579, -97.772880745, -97.77350612, -97.773500284, -97.807906757, 
    -97.8079127079999, -97.8085382949999, -97.808544248, -97.809169837, 
    -97.809175792, -97.809488587, -97.809494544, -97.80980734, 
    -97.8098132979999, -97.810126095, -97.810751689, -97.810763611, 
    -97.811389209, -97.811383246, -97.8120088429999, -97.812014807, 
    -97.812640405, -97.812646372, -97.813584772, -97.813590742, 
    -97.814216344, -97.814222316, -97.814535118, -97.814541091, 
    -97.814853894, -97.814859869, -97.815172672, -97.815178648, 
    -97.8154914529999, -97.8154974289999, -97.8167486519999, -97.816754633, 
    -97.817380246, -97.817386229, -97.818950267, -97.8189562539999, 
    -97.820520296, -97.820514303, -97.822703953, -97.822709953, 
    -97.826463646, -97.826457634, -97.8283344719999, -97.8283404909999, 
    -97.829278912, -97.829272891, -97.829898503, -97.829892479, 
    -97.830518089, -97.830512063, -97.831763278, -97.831769308, 
    -97.8327077229999, -97.832713756, -97.8330265609999, -97.833032596, 
    -97.833971016, -97.833977053, -97.8349154749999, -97.834921516, 
    -97.835859941, -97.8358659849999, -97.837430032, -97.83743608, 
    -97.838374511, -97.838380563, -97.8386933739999, -97.8386994269999, 
    -97.839950675, -97.839956733, -97.842146423, -97.842152487, 
    -97.8424653009999, -97.842477432, -97.842790248, -97.8427963139999, 
    -97.8431091309999, -97.843115199, -97.843428016, -97.843440154, 
    -97.843127334, -97.843145538, -97.842832715, -97.842850915, 
    -97.842538089, -97.842556287, -97.842243458, -97.8422677189999, 
    -97.841954885, -97.841973078, -97.8416602409999, -97.841678431, 
    -97.841365592, -97.841383779, -97.8410709359999, -97.8410769979999, 
    -97.8407641539999, -97.840770214, -97.841083059, -97.841089121, 
    -97.8407762749999, -97.840782335, -97.840469489, -97.840475548, 
    -97.8401627, -97.8401687589999, -97.83985591, -97.839861967, 
    -97.839549117, -97.83956123, -97.839248378, -97.839266545, -97.83895369, 
    -97.8389657989999, -97.838652942, -97.838658996, -97.838346137, 
    -97.83835219, -97.83803933, -97.838045382, -97.837732521, -97.837738572, 
    -97.83742571, -97.83743176, -97.836493172, -97.836499218, -97.83587349, 
    -97.8358795349999, -97.83494094, -97.834946982, -97.834008383, 
    -97.8340144209999, -97.833701554, -97.8337075919999, -97.833081855, 
    -97.8330878899999, -97.832775021, -97.832781056, -97.832468185, 
    -97.8324742189999, -97.832161347, -97.83216738, -97.8318545069999, 
    -97.831884666, -97.831571788, -97.831601942, -97.831289059, -97.83132524, 
    -97.831012351, -97.831157063, -97.830844149, -97.830850178, 
    -97.8305372629999, -97.830543291, -97.830230375, -97.830236402, 
    -97.829610567, -97.829616593, -97.829303674, -97.829309698, 
    -97.828996779, -97.829002802, -97.8286898809999, -97.828695904, 
    -97.8283829819999, -97.828389003, -97.8280760809999, -97.828082101, 
    -97.8277691769999, -97.8277751959999, -97.8274622709999, -97.82746829, 
    -97.827155364, -97.8271613809999, -97.826535527, -97.826541542, 
    -97.825915686, -97.825921699, -97.82560877, -97.8256147819999, 
    -97.8253018519999, -97.825307863, -97.824994932, -97.824682, 
    -97.824669982, -97.824357053, -97.824351045, -97.8240381159999, 
    -97.824032109, -97.823719182, -97.823713176, -97.82340025, -97.823394245, 
    -97.823081319, -97.823075316, -97.822762391, -97.8227563889999, 
    -97.822130542, -97.8221245409999, -97.821811619, -97.821805619, 
    -97.820866855, -97.8208608579999, -97.820235017, -97.820229023, 
    -97.819916103, -97.81991011, -97.818971354, -97.818965364, 
    -97.8180266109999, -97.818020624, -97.817081873, -97.817075889, 
    -97.816762973, -97.816756991, -97.816444076, -97.816432112, 
    -97.8161191999999, -97.816107238, -97.815794328, -97.815788348, 
    -97.815475438, -97.8154634809999, -97.815150574, -97.815144596, 
    -97.814831689, -97.8148197369999, -97.814506832, -97.814500857, 
    -97.814187953, -97.814181979, -97.8138690759999, -97.81385713, 
    -97.81354423, -97.8135382579999, -97.813225358, -97.8132193869999, 
    -97.812906488, -97.812900518, -97.812587621, -97.8125816519999, 
    -97.811955858, -97.811949892, -97.8116369959999, -97.8116310299999, 
    -97.811318135, -97.8113121709999, -97.810999277, -97.810993313, 
    -97.810680421, -97.8106744579999, -97.810361566, -97.810349644, 
    -97.809723864, -97.809717905, -97.809405016, -97.8093990579999, 
    -97.8090861699999, -97.809080213, -97.808767326, -97.80876137, 
    -97.8084484839999, -97.808442529, -97.808129644, -97.8081236899999, 
    -97.807810806, -97.807798901, -97.807486019, -97.807468165, 
    -97.807155286, -97.807119584, -97.806806711, -97.806794813, 
    -97.8064819419999, -97.806428411, -97.806115549, -97.806097709, 
    -97.8057848509999, -97.80577296, -97.805460103, -97.80544227, 
    -97.805129417, -97.8051115869999, -97.8054244369999, -97.805400661, 
    -97.805713507, -97.805701617, -97.806014461, -97.80597284, -97.805660003, 
    -97.8056243359999, -97.805311505, -97.805293675, -97.804980847, 
    -97.8049630199999, -97.805275845, -97.805246129, -97.805558949, 
    -97.8055292289999, -97.805216415, -97.805186701, -97.804873892, 
    -97.8048560669999, -97.804543261, -97.80452544, -97.8048382429999, 
    -97.8048263599999, -97.8051391609999, -97.805133219, -97.805446019, 
    -97.805440076, -97.805752874, -97.8057469299999, -97.806059728, 
    -97.806053783, -97.806366579, -97.8063606329999, -97.8066734289999, 
    -97.806667481, -97.8072930709999, -97.8072871209999, -97.807599915, 
    -97.807593964, -97.807906757, -97.852452724, -97.852458821, 
    -97.852146064, -97.852152161, -97.851839403, -97.851857689, 
    -97.851544928, -97.8515693049999, -97.85188207, -97.851894262, 
    -97.8522070289999, -97.852219222, -97.852531991, -97.852544187, 
    -97.852550285, -97.852237512, -97.852243609, -97.851618063, 
    -97.8516241569999, -97.8513113829999, -97.851317477, -97.851004701, 
    -97.851010794, -97.8506980179999, -97.850704109, -97.8500785539999, 
    -97.850084644, -97.849771865, -97.849777954, -97.849152394, 
    -97.849158481, -97.8475945759999, -97.847600658, -97.846975093, 
    -97.846981173, -97.846355606, -97.846361684, -97.846048899, 
    -97.846061053, -97.845748266, -97.845754342, -97.845441555, 
    -97.845447629, -97.8451348409999, -97.8451409149999, -97.844828125, 
    -97.84484027, -97.844527479, -97.844545694, -97.844232899, -97.844245041, 
    -97.843932244, -97.843956525, -97.843643723, -97.843661931, 
    -97.843349126, -97.843361263, -97.843048457, -97.843054524, 
    -97.842741716, -97.8427477829999, -97.842434974, -97.842447105, 
    -97.8421342939999, -97.842146423, -97.839956733, -97.839950675, 
    -97.8386994269999, -97.8386933739999, -97.838380563, -97.838374511, 
    -97.83743608, -97.837430032, -97.8358659849999, -97.835859941, 
    -97.834921516, -97.8349154749999, -97.833977053, -97.833971016, 
    -97.833032596, -97.8330265609999, -97.832713756, -97.8327077229999, 
    -97.831769308, -97.831763278, -97.830512063, -97.830518089, 
    -97.829892479, -97.829898503, -97.829272891, -97.829278912, 
    -97.8283404909999, -97.8283344719999, -97.826457634, -97.826463646, 
    -97.822709953, -97.822703953, -97.820514303, -97.820520296, 
    -97.8189562539999, -97.818950267, -97.817386229, -97.817380246, 
    -97.816754633, -97.8167486519999, -97.8154974289999, -97.8154914529999, 
    -97.815178648, -97.815172672, -97.814859869, -97.814853894, 
    -97.814541091, -97.814535118, -97.814222316, -97.814216344, 
    -97.813590742, -97.813584772, -97.812646372, -97.812640405, 
    -97.812014807, -97.8120088429999, -97.811383246, -97.811389209, 
    -97.810763611, -97.810751689, -97.810126095, -97.810120136, 
    -97.810432933, -97.8104210129999, -97.810733807, -97.810727847, 
    -97.812917397, -97.8129114289999, -97.813224221, -97.81323019, 
    -97.8169837, -97.8169896809999, -97.81886644, -97.818860452, 
    -97.82011162, -97.820105629, -97.82073121, -97.820725217, -97.821350796, 
    -97.821344801, -97.8219703779999, -97.8219643799999, -97.8238411039999, 
    -97.823835101, -97.824460673, -97.824454668, -97.8247674529999, 
    -97.824761446, -97.82507423, -97.825068222, -97.8253810049999, 
    -97.825374997, -97.825687779, -97.825681769, -97.829122356, 
    -97.829116335, -97.833495243, -97.833489207, -97.833801985, 
    -97.833795949, -97.834108726, -97.834102688, -97.8347282399999, 
    -97.8347222, -97.835034975, -97.835028935, -97.835341708, -97.835335667, 
    -97.835648439, -97.835642397, -97.8359551679999, -97.83626794, 
    -97.836261895, -97.836887436, -97.83688139, -97.837506928, 
    -97.8375008799999, -97.837813648, -97.837807598, -97.838120365, 
    -97.838114315, -97.838427081, -97.8384210299999, -97.838733794, 
    -97.8387277419999, -97.8390405059999, -97.839034453, -97.839659978, 
    -97.839653923, -97.840279446, -97.8402733889999, -97.840586149, 
    -97.8405800909999, -97.841831128, -97.841825066, -97.843076098, 
    -97.843070032, -97.8446338159999, -97.844627745, -97.846191523, 
    -97.846185447, -97.846498201, -97.846504279, -97.849944587, 
    -97.849938498, -97.8508767599999, -97.850882852, -97.851195607, 
    -97.8512017, -97.852452724, -97.8455203779999, -97.847083852, 
    -97.847089931, -97.847402626, -97.847408706, -97.847721403, 
    -97.847727483, -97.848040181, -97.8480523439999, -97.8486777429999, 
    -97.8486838269999, -97.848996528, -97.849002613, -97.8496280159999, 
    -97.849634103, -97.8499468049999, -97.849958981, -97.850271686, 
    -97.8502777749999, -97.850590481, -97.850596571, -97.850909277, 
    -97.8509153689999, -97.851228076, -97.851234169, -97.851546877, 
    -97.8515529699999, -97.8518656799999, -97.851871774, -97.853122616, 
    -97.853128715, -97.853441426, -97.8534353269999, -97.8537480369999, 
    -97.8537541379999, -97.854066849, -97.854072951, -97.854385663, 
    -97.854391766, -97.854704479, -97.854710583, -97.854397869, 
    -97.8544222799999, -97.854109562, -97.854121766, -97.853809045, 
    -97.85383345, -97.853520725, -97.853532925, -97.853220198, -97.853244595, 
    -97.853557326, -97.8536183319999, -97.853931073, -97.853973787, 
    -97.853661039, -97.85366714, -97.8533543899999, -97.85336659, 
    -97.853053839, -97.853066037, -97.852753283, -97.85276548, -97.852452724, 
    -97.8512017, -97.851195607, -97.850882852, -97.8508767599999, 
    -97.849938498, -97.849944587, -97.846504279, -97.846498201, 
    -97.846185447, -97.846191523, -97.844627745, -97.8446338159999, 
    -97.843070032, -97.843076098, -97.841825066, -97.841831128, 
    -97.8405800909999, -97.840586149, -97.8402733889999, -97.840279446, 
    -97.839653923, -97.839659978, -97.839034453, -97.8390405059999, 
    -97.8387277419999, -97.838733794, -97.8384210299999, -97.838427081, 
    -97.838114315, -97.838120365, -97.837807598, -97.837813648, 
    -97.8375008799999, -97.837506928, -97.83688139, -97.836887436, 
    -97.836261895, -97.83626794, -97.8359551679999, -97.835924953, 
    -97.835612187, -97.835606145, -97.8352933799999, -97.835287339, 
    -97.8346618099999, -97.834655771, -97.834343008, -97.834324895, 
    -97.8346376549999, -97.834631617, -97.834318857, -97.834300745, 
    -97.833987989, -97.83392159, -97.833909518, -97.834222261, 
    -97.8342101869999, -97.834522928, -97.83451689, -97.8348296299999, 
    -97.834823591, -97.8354490679999, -97.8354430269999, -97.8357557639999, 
    -97.83574368, -97.836369151, -97.836363107, -97.836675841, -97.836669796, 
    -97.836982529, -97.836970438, -97.837283169, -97.837277122, 
    -97.837589852, -97.837577757, -97.837890484, -97.837878387, 
    -97.8381911129999, -97.838185063, -97.838497788, -97.838491737, 
    -97.8388044609999, -97.838798409, -97.839111131, -97.839099026, 
    -97.839411747, -97.8394056929999, -97.839718412, -97.839712358, 
    -97.840025076, -97.840012965, -97.840325681, -97.840319625, -97.84125777, 
    -97.8412517099999, -97.841564424, -97.841558364, -97.841871077, 
    -97.841858954, -97.842171665, -97.84215954, -97.843410374, 
    -97.8434043079999, -97.843717015, -97.843710948, -97.844336361, 
    -97.8443302909999, -97.8446429969999, -97.844636926, -97.84494963, 
    -97.844931416, -97.8452441169999, -97.845238045, -97.845550745, 
    -97.8455203779999, -97.804347177, -97.804364985, -97.804677598, 
    -97.804683535, -97.804996149, -97.805002087, -97.805314702, 
    -97.805320641, -97.805633257, -97.8056391969999, -97.805951814, 
    -97.805963697, -97.806276315, -97.8062941429999, -97.806606765, 
    -97.806612709, -97.808488444, -97.808494394, -97.809432264, 
    -97.809438217, -97.811001339, -97.8110072969999, -97.811632547, 
    -97.811638508, -97.811951134, -97.811957095, -97.812582349, 
    -97.812588313, -97.8138388249999, -97.813832857, -97.814458111, 
    -97.814464081, -97.8147767089999, -97.814782679, -97.815407937, 
    -97.815401964, -97.81602722, -97.8160212449999, -97.816333871, 
    -97.816327895, -97.817265772, -97.817271751, -97.8175843769999, 
    -97.817590357, -97.818215612, -97.818221594, -97.818534223, 
    -97.818540206, -97.819165465, -97.8191714499999, -97.8194840799999, 
    -97.819490066, -97.819802698, -97.8198086849999, -97.820121317, 
    -97.820133294, -97.820758563, -97.8207525719999, -97.821065206, 
    -97.8210592139999, -97.821684478, -97.821678485, -97.825430055, 
    -97.8254360609999, -97.825748692, -97.825754699, -97.826067332, 
    -97.8260733399999, -97.826385973, -97.826397992, -97.826710627, 
    -97.8267166369999, -97.827029274, -97.827047308, -97.827359947, 
    -97.8273779849999, -97.827690627, -97.827696641, -97.828009285, 
    -97.828015299, -97.828327944, -97.82833396, -97.828646605, 
    -97.8286526219999, -97.828965269, -97.828971286, -97.829596582, 
    -97.829608621, -97.829921271, -97.829927292, -97.8305525929999, 
    -97.830558616, -97.830871268, -97.830877292, -97.8315025969999, 
    -97.831508623, -97.8321339299999, -97.832139959, -97.832765267, 
    -97.832771298, -97.833396608, -97.833402641, -97.834027954, 
    -97.8340400229999, -97.834352681, -97.834358717, -97.834671376, 
    -97.8346834499999, -97.834996111, -97.835002149, -97.835314812, 
    -97.8353329289999, -97.835645594, -97.8356576739999, -97.8359703419999, 
    -97.8359763829999, -97.8362890509999, -97.836301136, -97.8366138059999, 
    -97.83661985, -97.8369325209999, -97.836938566, -97.837251238, 
    -97.837257284, -97.837569957, -97.837588097, -97.8379007729999, 
    -97.837906821, -97.838219499, -97.8382376449999, -97.837924965, 
    -97.8379310129999, -97.8369929679999, -97.836999013, -97.8360609649999, 
    -97.8360670069999, -97.835128955, -97.835134994, -97.8348223089999, 
    -97.834828347, -97.833890289, -97.833896324, -97.832645575, 
    -97.832651606, -97.832338917, -97.832344947, -97.832032257, 
    -97.8320382859999, -97.831725596, -97.8317316229999, -97.831418932, 
    -97.8314249589999, -97.831112266, -97.831124318, -97.830811623, 
    -97.8308236729999, -97.830510976, -97.830517, -97.830204302, 
    -97.8302103249999, -97.829897626, -97.829909669, -97.829596968, 
    -97.82960901, -97.8292963069999, -97.8293083469999, -97.8289956419999, 
    -97.829001661, -97.828376248, -97.828382265, -97.8277568509999, 
    -97.8277628659999, -97.827450157, -97.8274561709999, -97.827143461, 
    -97.827149474, -97.826524053, -97.8265300639999, -97.825904641, 
    -97.82591065, -97.8255979369999, -97.825615961, -97.825303245, 
    -97.8253212659999, -97.825008547, -97.8250205589999, -97.8247078379999, 
    -97.824713843, -97.8244011209999, -97.8244071249999, -97.824094402, 
    -97.824100405, -97.8237876809999, -97.823793683, -97.8234809579999, 
    -97.823486959, -97.822861506, -97.822867505, -97.8213038659999, 
    -97.82130986, -97.820058945, -97.8200649349999, -97.819439474, 
    -97.819445462, -97.8178818059999, -97.8178877889999, -97.8175750569999, 
    -97.8175810389999, -97.817268305, -97.817274286, -97.816961552, 
    -97.816967532, -97.815716589, -97.815710613, -97.814146939, 
    -97.8141409679999, -97.8135154999999, -97.813503563, -97.813190831, 
    -97.8131848639999, -97.812246671, -97.812240706, -97.8119279759999, 
    -97.811922013, -97.811609284, -97.8116033219999, -97.811290594, 
    -97.811284632, -97.810971905, -97.810965945, -97.810653219, 
    -97.8106472599999, -97.810334535, -97.810322619, -97.8100098959999, 
    -97.810003939, -97.809691217, -97.809685261, -97.80937254, -97.809366586, 
    -97.8087411449999, -97.808735193, -97.8084224739999, -97.808416522, 
    -97.808103804, -97.8080978529999, -97.807785136, -97.8077791869999, 
    -97.8074664709999, -97.807460522, -97.806835092, -97.8068291449999, 
    -97.806516431, -97.806510486, -97.805885059, -97.805879116, 
    -97.805566404, -97.805560462, -97.805247751, -97.80524181, -97.804929099, 
    -97.80492316, -97.803985031, -97.803979095, -97.8030409689999, 
    -97.803035036, -97.802409621, -97.802403689, -97.8017782759999, 
    -97.801766417, -97.801453712, -97.8014418559999, -97.801129153, 
    -97.8011172989999, -97.800804598, -97.800798672, -97.800792746, 
    -97.801105445, -97.801099517, -97.801412215, -97.801406287, 
    -97.8017189829999, -97.8017130539999, -97.8020257489999, -97.802019819, 
    -97.8023325139999, -97.802326583, -97.802639276, -97.802633344, 
    -97.802946036, -97.802922304, -97.8032349919999, -97.8032231239999, 
    -97.802910438, -97.80289264, -97.802579957, -97.8025740259999, 
    -97.802261344, -97.802255413, -97.801942732, -97.801936803, 
    -97.801624123, -97.8016181949999, -97.801305516, -97.801293661, 
    -97.800980984, -97.8009750579999, -97.800349706, -97.800343782, 
    -97.8000311069999, -97.800025184, -97.7997125099999, -97.799706588, 
    -97.7990812419999, -97.799069402, -97.79844406, -97.7984381429999, 
    -97.798125473, -97.798119556, -97.7984322249999, -97.7984263069999, 
    -97.798738975, -97.7987330559999, -97.7990457229999, -97.799033884, 
    -97.7993465489999, -97.799305105, -97.798992447, -97.798974689, 
    -97.798662035, -97.798620608, -97.798307961, -97.798284294, 
    -97.798596937, -97.798537761, -97.7988503939999, -97.798826721, 
    -97.7985140919999, -97.79849634, -97.798808966, -97.798803048, 
    -97.799115672, -97.799080158, -97.799392777, -97.7993868569999, 
    -97.799699474, -97.7996935529999, -97.800318786, -97.800312863, 
    -97.800625478, -97.800619554, -97.800932168, -97.800926243, 
    -97.802489308, -97.802483378, -97.8027959899999, -97.802790059, 
    -97.803415281, -97.8034093479999, -97.804347177, -97.829836553, 
    -97.8301491349999, -97.8301551549999, -97.830467738, -97.830473759, 
    -97.8307863429999, -97.830792366, -97.831417535, -97.831423559, 
    -97.832048731, -97.832054757, -97.832367344, -97.832373372, 
    -97.832998547, -97.8330106069999, -97.833323196, -97.833329227, 
    -97.833954408, -97.833960441, -97.835210807, -97.8352168439999, 
    -97.8355294359999, -97.835535475, -97.835848068, -97.8358601469999, 
    -97.836172742, -97.8361848229999, -97.836497421, -97.836509504, 
    -97.836822103, -97.836840232, -97.836527629, -97.836539713, 
    -97.836227109, -97.836275437, -97.83658805, -97.836600134, -97.838475822, 
    -97.8384818709999, -97.839107102, -97.839113152, -97.839738385, 
    -97.839744438, -97.840057055, -97.840063109, -97.8419388189999, 
    -97.841932759, -97.842557993, -97.8425519309999, -97.842864548, 
    -97.842858485, -97.843483715, -97.84347765, -97.843790263, -97.843784198, 
    -97.8444094229999, -97.8444033549999, -97.844715967, -97.844709898, 
    -97.845022509, -97.845028579, -97.845653802, -97.845659874, 
    -97.8459724859999, -97.845990706, -97.8463033209999, -97.846321544, 
    -97.846634163, -97.8466463139999, -97.846958935, -97.846965011, 
    -97.848528119, -97.848534201, -97.848846823, -97.848852906, 
    -97.849790776, -97.8497968619999, -97.8507347349999, -97.850740824, 
    -97.851366075, -97.851372166, -97.851684792, -97.8516908839999, 
    -97.852003512, -97.8520156979999, -97.852328327, -97.852334422, 
    -97.852647052, -97.852695817, -97.852383178, -97.852389273, 
    -97.852076633, -97.852082727, -97.851770087, -97.851776179, 
    -97.851463538, -97.851469629, -97.851156987, -97.851169168, 
    -97.8508565229999, -97.8509052429999, -97.85059259, -97.850604768, 
    -97.850292113, -97.850298201, -97.849985545, -97.850015981, 
    -97.8497033199999, -97.849727666, -97.849415, -97.8494271709999, 
    -97.848489168, -97.84849525, -97.8481825819999, -97.848188663, 
    -97.847563323, -97.847569403, -97.846944061, -97.846950138, 
    -97.8466374659999, -97.8466496189999, -97.846336945, -97.846428082, 
    -97.846740771, -97.846759003, -97.8470716959999, -97.847083852, 
    -97.8455203779999, -97.8455143049999, -97.8452016109999, -97.845189467, 
    -97.844876775, -97.844864633, -97.8445519429999, -97.844539803, 
    -97.844227115, -97.844221047, -97.843595673, -97.843589606, 
    -97.8432769199999, -97.843264789, -97.8426394209999, -97.8426333579999, 
    -97.8423206749999, -97.8423146119999, -97.84200193, -97.841995869, 
    -97.841683188, -97.841677127, -97.841051767, -97.841045709, 
    -97.840107672, -97.840101617, -97.838850904, -97.838856955, 
    -97.8385442759999, -97.838550326, -97.8382376449999, -97.838219499, 
    -97.837906821, -97.8379007729999, -97.837588097, -97.837569957, 
    -97.837257284, -97.837251238, -97.836938566, -97.8369325209999, 
    -97.83661985, -97.8366138059999, -97.836301136, -97.8362890509999, 
    -97.8359763829999, -97.8359703419999, -97.8356576739999, -97.835645594, 
    -97.8353329289999, -97.835314812, -97.835002149, -97.834996111, 
    -97.8346834499999, -97.834671376, -97.834358717, -97.834352681, 
    -97.8340400229999, -97.834027954, -97.833402641, -97.833396608, 
    -97.832771298, -97.832765267, -97.832139959, -97.8321339299999, 
    -97.831508623, -97.8315025969999, -97.830877292, -97.830871268, 
    -97.830558616, -97.8305525929999, -97.829927292, -97.829921271, 
    -97.829608621, -97.829596582, -97.828971286, -97.828965269, 
    -97.8286526219999, -97.828646605, -97.82833396, -97.828327944, 
    -97.828015299, -97.828009285, -97.827696641, -97.827690627, 
    -97.8273779849999, -97.827359947, -97.827047308, -97.827029274, 
    -97.8267166369999, -97.826710627, -97.826397992, -97.826385973, 
    -97.8260733399999, -97.826067332, -97.825754699, -97.825748692, 
    -97.8254360609999, -97.825430055, -97.821678485, -97.821684478, 
    -97.8210592139999, -97.821065206, -97.8207525719999, -97.820758563, 
    -97.820133294, -97.820121317, -97.8198086849999, -97.819802698, 
    -97.819490066, -97.8194840799999, -97.8191714499999, -97.819165465, 
    -97.818540206, -97.818534223, -97.818221594, -97.818215612, 
    -97.817590357, -97.8175843769999, -97.817271751, -97.817265772, 
    -97.816327895, -97.816333871, -97.8160212449999, -97.81602722, 
    -97.815401964, -97.815407937, -97.814782679, -97.8147767089999, 
    -97.814464081, -97.814458111, -97.813832857, -97.8138388249999, 
    -97.812588313, -97.812582349, -97.811957095, -97.811951134, 
    -97.811638508, -97.811632547, -97.8110072969999, -97.811001339, 
    -97.809438217, -97.809432264, -97.808494394, -97.808488444, 
    -97.806612709, -97.806606765, -97.8062941429999, -97.806276315, 
    -97.805963697, -97.805951814, -97.8056391969999, -97.805633257, 
    -97.805320641, -97.805314702, -97.805002087, -97.804996149, 
    -97.804683535, -97.804677598, -97.804364985, -97.804347177, 
    -97.8046597859999, -97.804653849, -97.804966458, -97.80496052, 
    -97.805585734, -97.805579794, -97.8058924009999, -97.80588646, 
    -97.807762091, -97.8077561429999, -97.8093191629999, -97.809313211, 
    -97.809625813, -97.8096198599999, -97.810245063, -97.810239108, 
    -97.810864309, -97.810858352, -97.811170951, -97.8111590349999, 
    -97.811471632, -97.811459714, -97.811772309, -97.811754429, 
    -97.812067021, -97.812049137, -97.8123617259999, -97.812355764, 
    -97.813606116, -97.81360015, -97.8142253239999, -97.814219355, 
    -97.814531941, -97.814525972, -97.8151511409999, -97.815139199, 
    -97.815451782, -97.815439837, -97.815752418, -97.8157464449999, 
    -97.816059024, -97.8160530499999, -97.818866253, -97.81886027, 
    -97.8194854239999, -97.819491409, -97.8198039869999, -97.819809973, 
    -97.820435131, -97.8204471079999, -97.820759688, -97.820771668, 
    -97.822647164, -97.822641168, -97.8235789129999, -97.823572914, 
    -97.825135815, -97.825129811, -97.826380128, -97.8263861359999, 
    -97.826698716, -97.826710734, -97.827023316, -97.827035337, 
    -97.827660505, -97.827654492, -97.82952999, -97.829523971, -97.829836553, 
    -97.8354430269999, -97.8354490679999, -97.834823591, -97.8348296299999, 
    -97.83451689, -97.834522928, -97.8342101869999, -97.834222261, 
    -97.833909518, -97.83392159, -97.8336088459999, -97.833620916, 
    -97.833308169, -97.833314203, -97.833001455, -97.833025587, 
    -97.8327128349999, -97.8327249, -97.832412145, -97.832418177, 
    -97.8321054209999, -97.8321174819999, -97.832430239, -97.832472459, 
    -97.83184693, -97.83185296, -97.831540194, -97.831564309, -97.831877079, 
    -97.8318831079999, -97.832195879, -97.83220191, -97.832514682, 
    -97.8325207139999, -97.832833486, -97.8328395189999, -97.833152293, 
    -97.833158327, -97.833471102, -97.833477137, -97.833789913, 
    -97.833795949, -97.833801985, -97.833489207, -97.833495243, 
    -97.829116335, -97.829122356, -97.825681769, -97.82566975, -97.825356971, 
    -97.825332938, -97.825020163, -97.825014156, -97.8247013819999, 
    -97.824695376, -97.8243826029999, -97.824376598, -97.824063826, 
    -97.824057822, -97.8237450509999, -97.8237390479999, -97.823426279, 
    -97.823420277, -97.823107508, -97.823101507, -97.822788739, 
    -97.822782739, -97.8227767399999, -97.822463974, -97.822451977, 
    -97.823077504, -97.8230715029999, -97.8233842659999, -97.823378264, 
    -97.824003787, -97.823997784, -97.824310544, -97.82430454, -97.824617299, 
    -97.824611293, -97.826175085, -97.8261690739999, -97.827732859, 
    -97.8277268429999, -97.8283523549999, -97.828346337, -97.828659091, 
    -97.8286530729999, -97.8289658259999, -97.8289598059999, 
    -97.8295853119999, -97.82957929, -97.8298920409999, -97.829879996, 
    -97.830192745, -97.830186721, -97.8308122179999, -97.830806192, 
    -97.831118939, -97.831112912, -97.831425659, -97.831419631, 
    -97.831732376, -97.831726347, -97.832039091, -97.8320330609999, 
    -97.8323458039999, -97.832339774, -97.832652515, -97.832646484, 
    -97.832959224, -97.832953192, -97.833265932, -97.8332598979999, 
    -97.833572636, -97.833566602, -97.8354430269999, -97.83392159, 
    -97.833987989, -97.834300745, -97.834318857, -97.834631617, 
    -97.8346376549999, -97.834324895, -97.834343008, -97.834655771, 
    -97.8346618099999, -97.835287339, -97.8352933799999, -97.835606145, 
    -97.835612187, -97.835924953, -97.8359551679999, -97.835642397, 
    -97.835648439, -97.835335667, -97.835341708, -97.835028935, 
    -97.835034975, -97.8347222, -97.8347282399999, -97.834102688, 
    -97.834108726, -97.833795949, -97.833789913, -97.833477137, 
    -97.833471102, -97.833158327, -97.833152293, -97.8328395189999, 
    -97.832833486, -97.8325207139999, -97.832514682, -97.83220191, 
    -97.832195879, -97.8318831079999, -97.831877079, -97.831564309, 
    -97.831540194, -97.83185296, -97.83184693, -97.832472459, -97.832430239, 
    -97.8321174819999, -97.8321054209999, -97.832418177, -97.832412145, 
    -97.8327249, -97.8327128349999, -97.833025587, -97.833001455, 
    -97.833314203, -97.833308169, -97.833620916, -97.8336088459999, 
    -97.83392159, -97.798412537, -97.799037651, -97.7990435679999, 
    -97.799981241, -97.799987162, -97.800299721, -97.8003056429999, 
    -97.800618202, -97.800624125, -97.8009366859999, -97.8009426099999, 
    -97.801880295, -97.801874368, -97.802186928, -97.802192856, 
    -97.802505418, -97.802511347, -97.804074159, -97.804080093, 
    -97.8043926559999, -97.804398592, -97.8047111559999, -97.804717092, 
    -97.805967353, -97.805973294, -97.8062858599999, -97.806291802, 
    -97.8069169359999, -97.8069228799999, -97.807235448, -97.807241393, 
    -97.807553962, -97.807559908, -97.807872478, -97.807878425, 
    -97.810066421, -97.810691563, -97.810697519, -97.811010091, 
    -97.811022005, -97.8113345789999, -97.811340537, -97.812903411, 
    -97.812909374, -97.81322195, -97.813227915, -97.813540491, -97.813546457, 
    -97.8141716119999, -97.81417758, -97.814802737, -97.8148087069999, 
    -97.815121286, -97.815127257, -97.815439837, -97.815451782, 
    -97.815139199, -97.8151511409999, -97.814525972, -97.814531941, 
    -97.814219355, -97.8142253239999, -97.81360015, -97.813606116, 
    -97.812355764, -97.8123617259999, -97.812049137, -97.812067021, 
    -97.811754429, -97.811772309, -97.811459714, -97.811471632, 
    -97.8111590349999, -97.811170951, -97.810858352, -97.810864309, 
    -97.810239108, -97.810245063, -97.8096198599999, -97.809625813, 
    -97.809313211, -97.8093191629999, -97.8077561429999, -97.807762091, 
    -97.80588646, -97.8058924009999, -97.805579794, -97.805585734, 
    -97.80496052, -97.804966458, -97.804653849, -97.8046597859999, 
    -97.804347177, -97.8034093479999, -97.803415281, -97.802790059, 
    -97.8027959899999, -97.802483378, -97.802489308, -97.800926243, 
    -97.800932168, -97.800619554, -97.800625478, -97.800312863, 
    -97.800318786, -97.7996935529999, -97.799699474, -97.7993868569999, 
    -97.799392777, -97.799080158, -97.799115672, -97.798803048, 
    -97.798808966, -97.79849634, -97.7985140919999, -97.797263576, 
    -97.797257663, -97.796945035, -97.796903652, -97.79627841, -97.7962725, 
    -97.7959598799999, -97.795948063, -97.795635445, -97.79562363, 
    -97.795311014, -97.795299202, -97.794986588, -97.794957061, 
    -97.794644453, -97.794632645, -97.794320038, -97.794290523, 
    -97.793977922, -97.793960216, -97.793647618, -97.7936358169999, 
    -97.79332322, -97.793317321, -97.7930047249999, -97.792998827, 
    -97.7926862319999, -97.7926390539999, -97.7923264679999, 
    -97.7923146749999, -97.792002091, -97.7919903009999, -97.7916777189999, 
    -97.79164825, -97.791335673, -97.7913121019999, -97.790999529, 
    -97.790993638, -97.790368493, -97.7903626039999, -97.7900500329999, 
    -97.790044145, -97.789731574, -97.789725687, -97.789413118, 
    -97.789407232, -97.788782095, -97.788770327, -97.7890828929999, 
    -97.7890770079999, -97.789389574, -97.789383688, -97.7896962519999, 
    -97.789684478, -97.7899970399999, -97.789991152, -97.791866517, 
    -97.791860623, -97.794361099, -97.7943670019999, -97.795929803, 
    -97.795923896, -97.797174132, -97.7971682209999, -97.797793337, 
    -97.797787423, -97.798412537, -97.791624892, -97.791937411, 
    -97.791943304, -97.7922558239999, -97.792261718, -97.792574239, 
    -97.7925860299999, -97.792898553, -97.792916243, -97.7932287689999, 
    -97.793240565, -97.7932464629999, -97.793558992, -97.793564891, 
    -97.7938774199999, -97.79388332, -97.794195851, -97.794207654, 
    -97.7945201859999, -97.7945260879999, -97.794838622, -97.794844526, 
    -97.795469595, -97.795487311, -97.795174774, -97.795186583, 
    -97.795499122, -97.795505028, -97.795817569, -97.795864824, 
    -97.796177373, -97.796183281, -97.79680838, -97.7968202009999, 
    -97.797132753, -97.797138664, -97.7974512169999, -97.797457129, 
    -97.797769683, -97.797775596, -97.7980881509999, -97.798094066, 
    -97.798406621, -97.798412537, -97.797787423, -97.797793337, 
    -97.7971682209999, -97.797174132, -97.795923896, -97.795929803, 
    -97.7943670019999, -97.794361099, -97.791860623, -97.791866517, 
    -97.789991152, -97.788740908, -97.7887350239999, -97.788422464, 
    -97.788428346, -97.7881157849999, -97.788127549, -97.787502422, 
    -97.787508302, -97.786883173, -97.7868890509999, -97.785326223, 
    -97.785332096, -97.785019529, -97.785025401, -97.784712833, 
    -97.7847187039999, -97.784406135, -97.784423744, -97.7841111719999, 
    -97.78412291, -97.784128779, -97.7838162039999, -97.783822072, 
    -97.783509495, -97.7835153619999, -97.783202785, -97.7832086509999, 
    -97.782896073, -97.782901938, -97.7825893579999, -97.7825952219999, 
    -97.782282642, -97.782294368, -97.781981785, -97.781993509, 
    -97.781680925, -97.781686786, -97.7813742, -97.7813800599999, 
    -97.781067473, -97.78109091, -97.780778319, -97.7807958939999, 
    -97.7804833, -97.780489157, -97.780176562, -97.780170706, -97.779545517, 
    -97.779539663, -97.7789144769999, -97.778908625, -97.7779708479999, 
    -97.777976697, -97.776726324, -97.776732169, -97.776419574, 
    -97.776431262, -97.776118665, -97.7761303509999, -97.775817753, 
    -97.775829437, -97.775516836, -97.775522677, -97.775210075, 
    -97.775215915, -97.7742781059999, -97.7742722689999, -97.773334463, 
    -97.773328629, -97.772703427, -97.772697595, -97.772384995, 
    -97.772379164, -97.771441367, -97.771435539, -97.771122941, 
    -97.771111288, -97.770798692, -97.770792866, -97.7704802709999, 
    -97.770474447, -97.769536664, -97.769530843, -97.768905656, 
    -97.768899837, -97.7685872439999, -97.76856979, -97.76888238, 
    -97.7688591039999, -97.769171689, -97.76916005, -97.769472633, 
    -97.769431888, -97.769744464, -97.7697095349999, -97.7693969649999, 
    -97.769391145, -97.769078576, -97.7690727569999, -97.768760189, 
    -97.7687543709999, -97.768129238, -97.768123422, -97.767810856, 
    -97.767805041, -97.767492476, -97.767486662, -97.7671740979999, 
    -97.767168286, -97.766855723, -97.766849911, -97.766537349, 
    -97.766531538, -97.766519917, -97.766832476, -97.766815041, 
    -97.767127596, -97.767115971, -97.767428525, -97.7674227109999, 
    -97.767735264, -97.7677294489999, -97.768042001, -97.768036185, 
    -97.7686612859999, -97.768655468, -97.769593115, -97.769587295, 
    -97.770212391, -97.770206568, -97.770519115, -97.770513292, 
    -97.770825838, -97.770814189, -97.771126732, -97.7711150809999, 
    -97.771427623, -97.771410144, -97.771722682, -97.771716855, 
    -97.772029392, -97.7720235639999, -97.7723361, -97.772324442, 
    -97.7726369759999, -97.772631146, -97.772943679, -97.77294951, 
    -97.773574579, -97.7735804119999, -97.774518018, -97.774512181, 
    -97.774824715, -97.774830553, -97.7751430879999, -97.775148927, 
    -97.775773999, -97.7757798389999, -97.776404913, -97.776410756, 
    -97.777035832, -97.7770416769999, -97.777354216, -97.777360062, 
    -97.7776726019999, -97.777678449, -97.77830353, -97.778309379, 
    -97.779872088, -97.7798662339999, -97.780178774, -97.7801729189999, 
    -97.780485459, -97.7804796029999, -97.7807921409999, -97.780786284, 
    -97.7829740449999, -97.7829681809999, -97.783593253, -97.783587386, 
    -97.784524991, -97.7845191219999, -97.7848316559999, -97.784825785, 
    -97.785450851, -97.785444978, -97.788570294, -97.788564411, 
    -97.788876941, -97.7888710569999, -97.789183587, -97.789177702, 
    -97.78949023, -97.789478459, -97.789790985, -97.789785098, -97.790097623, 
    -97.790091736, -97.7904042599999, -97.790398371, -97.790710894, 
    -97.790705005, -97.791017526, -97.791011636, -97.791324157, 
    -97.791312374, -97.791624892 ;

 catchments_y = 30.3943565530001, 30.395706825, 30.3957120690001, 
    30.3959821230001, 30.395987367, 30.396797528, 30.3968027710001, 
    30.3970728240001, 30.3970780660001, 30.3973481190001, 30.3973586010001, 
    30.3976286540001, 30.397633893, 30.397903946, 30.3979248950001, 
    30.398465, 30.398470235, 30.3990103400001, 30.399015574, 
    30.3992856260001, 30.3992908600001, 30.399560912, 30.399576606, 
    30.3998466580001, 30.3998518880001, 30.400391991, 30.4003972200001, 
    30.4006672720001, 30.4006725, 30.4009425510001, 30.400947778, 
    30.40148788, 30.4014931070001, 30.4017631570001, 30.401768383, 
    30.4020384340001, 30.402043658, 30.4023137090001, 30.4023189320001, 
    30.402859033, 30.402864256, 30.4034043560001, 30.403409578, 
    30.4036796280001, 30.4036848490001, 30.404224948, 30.404230168, 
    30.4045002180001, 30.4045054370001, 30.4047754860001, 30.404785922, 
    30.4053260200001, 30.405331237, 30.4053625190001, 30.405632568, 
    30.405637778, 30.4059078270001, 30.4059130370001, 30.4061830850001, 
    30.4061882940001, 30.4064583430001, 30.4064635510001, 30.4067335990001, 
    30.4067388060001, 30.407008854, 30.4070140600001, 30.4072841080001, 
    30.407289314, 30.407559361, 30.4075645660001, 30.407834614, 30.407839817, 
    30.408109865, 30.4081202690001, 30.4083903170001, 30.4083955180001, 
    30.4089356120001, 30.408940812, 30.409210859, 30.4092212570001, 
    30.409491303, 30.409496501, 30.4097665480001, 30.4097717440001, 
    30.410041791, 30.410052181, 30.410322228, 30.4103481880001, 
    30.4106182350001, 30.410644173, 30.4109142190001, 30.410919404, 
    30.4111894500001, 30.4111946350001, 30.411464681, 30.4114750460001, 
    30.411745092, 30.411750274, 30.4120203200001, 30.41203068, 30.412570771, 
    30.412565591, 30.4128356370001, 30.4128459950001, 30.4125759500001, 
    30.4125966570001, 30.412326611, 30.412331785, 30.4112516020001, 
    30.411256775, 30.410716682, 30.4107218550001, 30.4104518080001, 
    30.41045698, 30.410186933, 30.410192104, 30.4099220570001, 30.409927226, 
    30.4096571790001, 30.409662348, 30.4077720130001, 30.407777181, 
    30.407237084, 30.4072422510001, 30.4069722020001, 30.4069773690001, 
    30.4053570720001, 30.4053622380001, 30.4045520870001, 30.404557251, 
    30.404287201, 30.404282037, 30.4040119860001, 30.4040068210001, 
    30.40373677, 30.403731604, 30.403461554, 30.4034357100001, 
    30.4031656600001, 30.403155316, 30.4028852650001, 30.4028645670001, 
    30.4025945160001, 30.402568624, 30.4022985730001, 30.4022882100001, 
    30.4020181590001, 30.402012976, 30.4017429250001, 30.401737741, 
    30.4014676890001, 30.401462505, 30.4011924530001, 30.4011872670001, 
    30.400917216, 30.400912029, 30.4003719250001, 30.4003667380001, 
    30.39955658, 30.399551392, 30.3987412330001, 30.398736044, 30.398465991, 
    30.398455611, 30.398185557, 30.398175173, 30.3979051200001, 30.397899927, 
    30.397629873, 30.397624679, 30.397354625, 30.3973442340001, 
    30.3970741800001, 30.397063786, 30.3967937310001, 30.3967885330001, 
    30.3962484240001, 30.396243225, 30.3957031160001, 30.395697915, 
    30.395157806, 30.395152604, 30.394882549, 30.394877347, 30.394607292, 
    30.394602089, 30.394061978, 30.394056774, 30.3935166630001, 30.393511458, 
    30.3932414020001, 30.3932361970001, 30.392966141, 30.392960934, 
    30.3926908780001, 30.392685671, 30.3924156140001, 30.3924104060001, 
    30.39214035, 30.3921195080001, 30.391849452, 30.3918338120001, 
    30.3915637550001, 30.3915585400001, 30.391288483, 30.391272832, 
    30.3910027750001, 30.3909871160001, 30.3907170590001, 30.390701393, 
    30.3904313350001, 30.3904261110001, 30.3904208860001, 30.390150829, 
    30.3901456030001, 30.389875546, 30.3898546340001, 30.390124691, 
    30.3901089980001, 30.390379056, 30.390368589, 30.3906386460001, 
    30.3906334120001, 30.3909034690001, 30.390898233, 30.3911682900001, 
    30.3911630530001, 30.39143311, 30.391422634, 30.391962747, 
    30.3919575080001, 30.3922275640001, 30.392217083, 30.392487139, 
    30.392481897, 30.393022009, 30.3930167660001, 30.393556877, 
    30.3935516330001, 30.394091743, 30.394086498, 30.3943565530001, 
    30.3582615230001, 30.358531602, 30.3585366890001, 30.3590768460001, 
    30.359081932, 30.3593520100001, 30.3593570960001, 30.359627174, 
    30.359632258, 30.359637342, 30.3599074200001, 30.3599175850001, 
    30.360187663, 30.3601927440001, 30.3604628210001, 30.3604780590001, 
    30.360748137, 30.3607735160001, 30.361043593, 30.361048666, 
    30.3613187440001, 30.361323816, 30.3615938930001, 30.3615989640001, 
    30.36105881, 30.3610537390001, 30.3602435060001, 30.3602384340001, 
    30.359968356, 30.3599632830001, 30.3596932040001, 30.3596881300001, 
    30.359418052, 30.359392669, 30.3591225910001, 30.3591124320001, 
    30.3588423530001, 30.35883219, 30.3582920330001, 30.35828695, 
    30.3580168710001, 30.3580117880001, 30.358281866, 30.3582615230001, 
    30.373633951, 30.373904021, 30.3738939290001, 30.374164, 
    30.3741589530001, 30.3744290230001, 30.3744239750001, 30.3746940450001, 
    30.374688996, 30.374959066, 30.374933807, 30.375203877, 30.3751988230001, 
    30.3754688920001, 30.375463837, 30.3757339060001, 30.37572885, 
    30.375998919, 30.375993862, 30.376263931, 30.3762487550001, 30.376518823, 
    30.376508701, 30.3762386330001, 30.3762234430001, 30.375413236, 
    30.3754081710001, 30.3751381020001, 30.3751330360001, 30.375403105, 
    30.375347322, 30.375617391, 30.3756123150001, 30.375882383, 
    30.3758722270001, 30.3761422960001, 30.3761372170001, 30.376407285, 
    30.376402205, 30.3766722730001, 30.3766671920001, 30.37693726, 
    30.3769321780001, 30.377202246, 30.3771971630001, 30.377467231, 
    30.3774112610001, 30.3771411930001, 30.3771361, 30.3768660320001, 
    30.3768609380001, 30.37659087, 30.376585775, 30.3763157070001, 
    30.3763106110001, 30.376040543, 30.3760252490001, 30.375755181, 
    30.3757296740001, 30.375999742, 30.3759895330001, 30.3762596010001, 
    30.3762544950001, 30.375984427, 30.3759793200001, 30.3759742120001, 
    30.37624428, 30.3762238410001, 30.3762187290001, 30.3772989980001, 
    30.3773041110001, 30.380004775, 30.380009886, 30.3810901470001, 
    30.3810850360001, 30.3829754870001, 30.382970374, 30.3837805650001, 
    30.3837754520001, 30.385665891, 30.3856710050001, 30.3862111290001, 
    30.386216242, 30.3864863040001, 30.386491415, 30.3867614770001, 
    30.3867665880001, 30.38703665, 30.3870315390001, 30.3873016000001, 
    30.3872913760001, 30.387831498, 30.3878212700001, 30.3880913310001, 
    30.388086216, 30.388356276, 30.3883511600001, 30.3886212210001, 
    30.3886109850001, 30.3888810460001, 30.3888759270001, 30.3894160470001, 
    30.389410927, 30.3896809870001, 30.3896758660001, 30.3899459260001, 
    30.389940804, 30.390210864, 30.390205741, 30.3904758, 30.3904706770001, 
    30.3912808540001, 30.3912757300001, 30.391815847, 30.3918209710001, 
    30.3929012040001, 30.392906328, 30.3931763860001, 30.3931815080001, 
    30.3934515660001, 30.3934566880001, 30.393726745, 30.3937318660001, 
    30.3940019240001, 30.394007044, 30.3942771010001, 30.394282221, 
    30.394552278, 30.394557396, 30.3948274530001, 30.3948581450001, 
    30.394588088, 30.394603422, 30.394333364, 30.394343582, 30.3940735250001, 
    30.394078633, 30.393808575, 30.393818788, 30.3935487300001, 
    30.3935742460001, 30.3933041880001, 30.393319487, 30.3935895450001, 
    30.3935997400001, 30.393869798, 30.393885084, 30.3936150260001, 
    30.393620119, 30.393350061, 30.3933551540001, 30.3930850950001, 
    30.393095278, 30.392825219, 30.392835398, 30.39256534, 30.392575515, 
    30.392305456, 30.3923105420001, 30.3917704240001, 30.3917755090001, 
    30.390695271, 30.390700355, 30.3890799930001, 30.3890850770001, 
    30.388815016, 30.38882518, 30.388555119, 30.388560199, 30.3882901380001, 
    30.3882952180001, 30.3880251570001, 30.388035314, 30.3877652520001, 
    30.3877804810001, 30.3872403570001, 30.3872454310001, 30.386975369, 
    30.386985515, 30.3867154530001, 30.386720525, 30.386450462, 30.386460603, 
    30.38619054, 30.386231068, 30.3859610050001, 30.385966067, 
    30.3856960040001, 30.3857415210001, 30.385776874, 30.385506811, 
    30.3855169030001, 30.38524684, 30.3852518850001, 30.3849818210001, 
    30.3849919080001, 30.3847218440001, 30.3847268860001, 30.3844568220001, 
    30.3844618640001, 30.3841917990001, 30.3841968400001, 30.3839267750001, 
    30.383931815, 30.38366175, 30.3836818990001, 30.3834118350001, 
    30.383421904, 30.3831518390001, 30.3831619050001, 30.382621774, 
    30.382626805, 30.38235674, 30.38236177, 30.3818216380001, 30.381826668, 
    30.3812865360001, 30.381291565, 30.3810214980001, 30.381026526, 
    30.3807564590001, 30.3807514310001, 30.380481365, 30.3804713060001, 
    30.3799311720001, 30.379926142, 30.379656074, 30.379651043, 
    30.3788408400001, 30.3788358080001, 30.3780256040001, 30.378020571, 
    30.3774804340001, 30.3774754, 30.3766651940001, 30.376660159, 
    30.3758499510001, 30.3758449160001, 30.3755748460001, 30.3755698100001, 
    30.3752997400001, 30.3752947020001, 30.3750246330001, 30.375019594, 
    30.374749524, 30.3747444850001, 30.3744744150001, 30.374469375, 
    30.374199305, 30.374189222, 30.373919152, 30.3739090660001, 
    30.3736389950001, 30.373633951, 30.359632258, 30.360172414, 30.360162244, 
    30.3604323210001, 30.360427235, 30.3606973120001, 30.360692225, 
    30.3609623020001, 30.3609572140001, 30.361227291, 30.3612171120001, 
    30.3614871890001, 30.3614820980001, 30.3625624040001, 30.362557312, 
    30.3639076910001, 30.363902598, 30.364442748, 30.364437654, 30.364977804, 
    30.3649727100001, 30.3671333020001, 30.3671282060001, 30.36739828, 
    30.367393183, 30.3676632560001, 30.367658159, 30.368198304, 
    30.3681932060001, 30.369003424, 30.3689983240001, 30.370348683, 
    30.3703435830001, 30.370883726, 30.370878625, 30.3722289780001, 
    30.3722238760001, 30.3727640160001, 30.372758913, 30.373299053, 
    30.3732939490001, 30.373834088, 30.3738289830001, 30.3740990520001, 
    30.3740888400001, 30.3759793200001, 30.375984427, 30.3762544950001, 
    30.3762596010001, 30.3759895330001, 30.375999742, 30.3757296740001, 
    30.375755181, 30.3760252490001, 30.376040543, 30.3763106110001, 
    30.3763157070001, 30.376585775, 30.37659087, 30.3768609380001, 
    30.3768660320001, 30.3771361, 30.3771411930001, 30.3774112610001, 
    30.377467231, 30.3771971630001, 30.377202246, 30.3769321780001, 
    30.37693726, 30.3766671920001, 30.3766722730001, 30.376402205, 
    30.376407285, 30.3761372170001, 30.3761422960001, 30.3758722270001, 
    30.375882383, 30.3756123150001, 30.375617391, 30.375347322, 30.375403105, 
    30.3751330360001, 30.3751381020001, 30.3754081710001, 30.375413236, 
    30.3762234430001, 30.3762386330001, 30.376508701, 30.376518823, 
    30.3762487550001, 30.376263931, 30.375993862, 30.375998919, 30.37572885, 
    30.3757339060001, 30.375463837, 30.3754688920001, 30.3751988230001, 
    30.375203877, 30.374933807, 30.374959066, 30.374688996, 30.3746940450001, 
    30.3744239750001, 30.3744290230001, 30.3741589530001, 30.374164, 
    30.3738939290001, 30.373904021, 30.373633951, 30.3728237380001, 
    30.372828783, 30.3714784250001, 30.371473381, 30.369852947, 
    30.3698479020001, 30.369037683, 30.3687676100001, 30.3687625640001, 
    30.3684924900001, 30.368487443, 30.3679472960001, 30.3679422480001, 
    30.3674021, 30.3673970520001, 30.366856903, 30.3668518540001, 
    30.3665817790001, 30.3665615730001, 30.3662914980001, 30.3662763340001, 
    30.366546408, 30.3665362950001, 30.3668063690001, 30.366796251, 
    30.367066326, 30.3670612650001, 30.3667911910001, 30.36678613, 
    30.3659759070001, 30.365970845, 30.364890545, 30.364885482, 30.364615407, 
    30.364610343, 30.364340268, 30.3643352030001, 30.3637950520001, 
    30.3637899870001, 30.363249834, 30.3632447680001, 30.362974692, 
    30.3629696250001, 30.362699548, 30.3626944810001, 30.362424404, 
    30.362419335, 30.362149259, 30.362144189, 30.3618741120001, 30.361869042, 
    30.3615989640001, 30.3615938930001, 30.361323816, 30.3613187440001, 
    30.361048666, 30.361043593, 30.3607735160001, 30.360748137, 
    30.3604780590001, 30.3604628210001, 30.3601927440001, 30.360187663, 
    30.3599175850001, 30.3599074200001, 30.359637342, 30.359632258, 
    30.382626805, 30.382631836, 30.38236177, 30.38235674, 30.382626805, 
    30.382626805, 30.382621774, 30.3831619050001, 30.3831518390001, 
    30.383421904, 30.3834118350001, 30.3836818990001, 30.38366175, 
    30.383931815, 30.3839267750001, 30.3841968400001, 30.3841917990001, 
    30.3844618640001, 30.3844568220001, 30.3847268860001, 30.3847218440001, 
    30.3849919080001, 30.3849818210001, 30.3852518850001, 30.38524684, 
    30.3855169030001, 30.385506811, 30.385776874, 30.3857415210001, 
    30.3860115850001, 30.3860469370001, 30.3863170010001, 30.3863220480001, 
    30.386592111, 30.386597157, 30.3876774070001, 30.387682453, 
    30.3879525150001, 30.387957559, 30.3882276210001, 30.388232665, 
    30.3885027270001, 30.3885077690001, 30.388777831, 30.388782873, 
    30.390673302, 30.390678343, 30.390948403, 30.3912184640001, 
    30.3912285430001, 30.3914986030001, 30.391503642, 30.391773702, 
    30.3917837760001, 30.3920538360001, 30.3920588710001, 30.3923289310001, 
    30.392333966, 30.3926040260001, 30.3926191250001, 30.3928891840001, 
    30.3928992460001, 30.392359126, 30.392364156, 30.390473732, 
    30.3904787600001, 30.390208699, 30.3902137270001, 30.389943665, 
    30.3899486920001, 30.389138507, 30.3891334800001, 30.386702917, 
    30.3866978900001, 30.386157763, 30.3861527350001, 30.384802415, 
    30.3847973860001, 30.3839871920001, 30.3839821620001, 30.3829019020001, 
    30.3828968710001, 30.382626805, 30.4157631570001, 30.4160332010001, 
    30.416038342, 30.416308386, 30.4163135260001, 30.417393701, 30.41739884, 
    30.417938926, 30.417944065, 30.4192942780001, 30.4192994150001, 
    30.4195694580001, 30.419574594, 30.4198446360001, 30.4198549070001, 
    30.4201249490001, 30.4201300830001, 30.4204001250001, 30.4204052580001, 
    30.420675299, 30.4206804310001, 30.4209504730001, 30.420955604, 
    30.420145479, 30.4201403480001, 30.4193302210001, 30.419325089, 
    30.419055047, 30.419049914, 30.4179697430001, 30.417964609, 30.417154479, 
    30.4171493440001, 30.416069168, 30.4160640330001, 30.4157939890001, 
    30.4157631570001, 30.3857415210001, 30.3856960040001, 30.385966067, 
    30.3859610050001, 30.386231068, 30.38619054, 30.386460603, 30.386450462, 
    30.386720525, 30.3867154530001, 30.386985515, 30.386975369, 
    30.3872454310001, 30.3872403570001, 30.3877804810001, 30.3877652520001, 
    30.388035314, 30.3880251570001, 30.3882952180001, 30.3882901380001, 
    30.388560199, 30.388555119, 30.38882518, 30.388815016, 30.3890850770001, 
    30.3890799930001, 30.390700355, 30.390695271, 30.3917755090001, 
    30.3917704240001, 30.3923105420001, 30.392305456, 30.392575515, 
    30.39256534, 30.392835398, 30.392825219, 30.393095278, 30.3930850950001, 
    30.3933551540001, 30.393350061, 30.393620119, 30.3936150260001, 
    30.393885084, 30.393869798, 30.3935997400001, 30.3935895450001, 
    30.393319487, 30.3933041880001, 30.3935742460001, 30.3935487300001, 
    30.393818788, 30.393808575, 30.394078633, 30.3940735250001, 30.394343582, 
    30.394333364, 30.394603422, 30.394588088, 30.3948581450001, 
    30.3948274530001, 30.39509751, 30.395092391, 30.395632504, 
    30.3956273850001, 30.3961674970001, 30.3961623770001, 30.3967024890001, 
    30.396692246, 30.396962301, 30.396952055, 30.39722211, 30.3972067330001, 
    30.3974767880001, 30.3974614030001, 30.3977314580001, 30.397726328, 
    30.3979963830001, 30.3979912520001, 30.398261307, 30.398256175, 
    30.398526229, 30.3985159630001, 30.3987860170001, 30.398780883, 
    30.399050937, 30.399040665, 30.399310719, 30.3993055820001, 
    30.3995756350001, 30.3995704970001, 30.3998405510001, 30.3998354120001, 
    30.400105465, 30.400100325, 30.400370378, 30.400360096, 30.4006301490001, 
    30.400625006, 30.4008950590001, 30.4008899150001, 30.4011599680001, 
    30.4011548240001, 30.401694929, 30.4016897830001, 30.4019598360001, 
    30.401954689, 30.4022247410001, 30.402219594, 30.402489646, 30.402484498, 
    30.4027545500001, 30.4027494010001, 30.403019452, 30.403014302, 
    30.4032843540001, 30.4032688990001, 30.40353895, 30.403533796, 
    30.404073898, 30.404063588, 30.4043336390001, 30.4043078490001, 
    30.4045779, 30.404557251, 30.4045520870001, 30.4053622380001, 
    30.4053570720001, 30.4069773690001, 30.4069722020001, 30.4072422510001, 
    30.407237084, 30.407777181, 30.4077720130001, 30.409662348, 
    30.4096675160001, 30.410207611, 30.4102179440001, 30.410758038, 
    30.410763203, 30.411573343, 30.4115785070001, 30.4118485540001, 
    30.411874363, 30.4121444090001, 30.412154727, 30.4124247730001, 
    30.4124299310001, 30.412699977, 30.4127154440001, 30.41298549, 
    30.412990644, 30.4135307350001, 30.41354104, 30.4138110850001, 
    30.413826537, 30.414366627, 30.4143717760001, 30.4149118650001, 
    30.414927306, 30.4151973510001, 30.4152024960001, 30.4152127840001, 
    30.4154828280001, 30.4154879710001, 30.4157580150001, 30.4157631570001, 
    30.4157939890001, 30.4160640330001, 30.416069168, 30.4171493440001, 
    30.417154479, 30.417964609, 30.4179697430001, 30.419049914, 30.419055047, 
    30.419325089, 30.4193302210001, 30.4201403480001, 30.420145479, 
    30.420955604, 30.421225646, 30.4212307760001, 30.421500817, 
    30.4215059470001, 30.4220460290001, 30.422051158, 30.4228612800001, 
    30.4228561510001, 30.4236662710001, 30.4236611420001, 30.425011339, 
    30.4250062090001, 30.4263564020001, 30.426361533, 30.4277117230001, 
    30.427716853, 30.4285269650001, 30.428521835, 30.4293319450001, 
    30.429326814, 30.4309470310001, 30.4309418990001, 30.4328321450001, 
    30.432837277, 30.433377346, 30.4333824770001, 30.4344626130001, 
    30.434467743, 30.4352778430001, 30.4352727130001, 30.4360828120001, 
    30.436077681, 30.436617746, 30.4366126140001, 30.4374227100001, 
    30.4374175770001, 30.4398478580001, 30.439842723, 30.4403827840001, 
    30.440377649, 30.4419978270001, 30.4419926910001, 30.442802778, 
    30.442797641, 30.4433376980001, 30.44333256, 30.4436025890001, 
    30.44359745, 30.4438674780001, 30.4438623390001, 30.4441323660001, 
    30.444127226, 30.444397254, 30.4443921120001, 30.44466214, 30.444656998, 
    30.444927025, 30.4449167380001, 30.4454567920001, 30.445451647, 
    30.445721674, 30.445716528, 30.445986555, 30.4459814080001, 
    30.4462514350001, 30.4462462870001, 30.4465163130001, 30.4465111650001, 
    30.4467811910001, 30.446770891, 30.447040917, 30.447087239, 
    30.4473572650001, 30.447367549, 30.447097523, 30.447112942, 
    30.4473829680001, 30.4474035150001, 30.447673541, 30.4476838090001, 
    30.4474137830001, 30.4474240480001, 30.447694074, 30.447724846, 
    30.447994872, 30.4480307320001, 30.4477607060001, 30.4477709440001, 
    30.4475009180001, 30.4475316100001, 30.4472615830001, 30.447292243, 
    30.44756227, 30.447592898, 30.447322871, 30.447338173, 30.447068146, 
    30.447078343, 30.446808316, 30.446823604, 30.446553577, 30.446558671, 
    30.446288644, 30.44629883, 30.4460288020001, 30.446033894, 
    30.4457638660001, 30.445774047, 30.4455040190001, 30.4455091080001, 
    30.4452390800001, 30.445244168, 30.4449741400001, 30.4449843130001, 
    30.444714285, 30.44471937, 30.444449342, 30.4444595100001, 30.444189481, 
    30.4441945630001, 30.4439245340001, 30.443929616, 30.442849499, 
    30.442854579, 30.441774459, 30.441779539, 30.4412394780001, 
    30.4412445570001, 30.440974526, 30.4409796040001, 30.440439542, 
    30.4404446190001, 30.440174588, 30.440179664, 30.4396396010001, 
    30.439644677, 30.439374645, 30.439379719, 30.438839655, 30.438844729, 
    30.438574697, 30.4385797690001, 30.4383097370001, 30.438314808, 
    30.438044776, 30.4380498470001, 30.4377798140001, 30.4377950210001, 
    30.4375249880001, 30.437530055, 30.4378000880001, 30.4378102200001, 
    30.437540187, 30.4375452520001, 30.4378152850001, 30.4378254110001, 
    30.4380954440001, 30.4381005060001, 30.4383705390001, 30.4383806600001, 
    30.4386506930001, 30.438655752, 30.438925785, 30.4389359, 30.439205933, 
    30.4392211000001, 30.4389510680001, 30.438956122, 30.438686089, 
    30.438696194, 30.438426162, 30.4384312130001, 30.4381611800001, 
    30.43816623, 30.4381712800001, 30.4379012470001, 30.4379062950001, 
    30.4376362620001, 30.4376413100001, 30.4373712760001, 30.437381369, 
    30.4371113350001, 30.4371214240001, 30.4368513910001, 30.436856434, 
    30.4365864000001, 30.4365964830001, 30.436326449, 30.43633149, 
    30.4360614550001, 30.4360715340001, 30.435801499, 30.4358115740001, 
    30.435541539, 30.435546575, 30.4352765400001, 30.43528661, 
    30.4350165750001, 30.43502664, 30.4347566050001, 30.4347616370001, 
    30.434491601, 30.4345016620001, 30.434231626, 30.434241683, 
    30.4339716470001, 30.4339766740001, 30.433706638, 30.4337166890001, 
    30.433446653, 30.4334567010001, 30.4331866650001, 30.433191687, 
    30.4329216510001, 30.4329316930001, 30.432661657, 30.432121583, 
    30.432116562, 30.4315764880001, 30.431571466, 30.431301429, 
    30.4312964060001, 30.4310263680001, 30.431021345, 30.430751307, 
    30.4307462830001, 30.430206207, 30.4302011820001, 30.4299311440001, 
    30.429926118, 30.42965608, 30.429651053, 30.429381015, 30.4293759870001, 
    30.428835909, 30.4288308810001, 30.4280207640001, 30.428015734, 
    30.4277456950001, 30.427740665, 30.4274706250001, 30.4274655940001, 
    30.4269255150001, 30.4269204830001, 30.426650443, 30.42664541, 
    30.4263753700001, 30.426370336, 30.4261002960001, 30.4260952610001, 
    30.425825221, 30.4258201850001, 30.425550145, 30.4255451080001, 
    30.4252750680001, 30.4252599530001, 30.4249899120001, 30.424984872, 
    30.4247148310001, 30.4247097910001, 30.42443975, 30.4244044390001, 
    30.424134398, 30.4241040970001, 30.423834056, 30.423829003, 
    30.4235589620001, 30.4235488530001, 30.42300877, 30.4230037140001, 
    30.422193588, 30.4221885310001, 30.420838319, 30.420833261, 30.420023132, 
    30.4200180730001, 30.4194779860001, 30.4194830450001, 30.418402869, 
    30.41839781, 30.4178577210001, 30.417852662, 30.417042528, 
    30.4170475870001, 30.416777542, 30.4167826, 30.4165125540001, 
    30.4165176120001, 30.416247566, 30.416242509, 30.415702418, 30.415697359, 
    30.41326694, 30.413271998, 30.4130019510001, 30.4130070080001, 
    30.4127369600001, 30.412742017, 30.412471969, 30.4124770240001, 
    30.411936928, 30.4119419830001, 30.411671934, 30.4116820400001, 
    30.4114119920001, 30.4114170440001, 30.411146995, 30.411152046, 
    30.4103418990001, 30.410336849, 30.4087165510001, 30.4087216020001, 
    30.4081815010001, 30.408186551, 30.407376399, 30.407381448, 
    30.4054910880001, 30.4054961360001, 30.403065661, 30.403060613, 
    30.40144029, 30.401445338, 30.400095064, 30.400100111, 30.3992899450001, 
    30.39929499, 30.397404597, 30.3974096420001, 30.3944390080001, 
    30.394433963, 30.393893846, 30.3938888010001, 30.3930786240001, 
    30.3930735770001, 30.3917232790001, 30.3917283260001, 30.391458265, 
    30.3914633110001, 30.3911932500001, 30.3912134230001, 30.390943362, 
    30.390948403, 30.390678343, 30.390673302, 30.388782873, 30.388777831, 
    30.3885077690001, 30.3885027270001, 30.388232665, 30.3882276210001, 
    30.387957559, 30.3879525150001, 30.387682453, 30.3876774070001, 
    30.386597157, 30.386592111, 30.3863220480001, 30.3863170010001, 
    30.3860469370001, 30.3860115850001, 30.3857415210001, 30.4152024960001, 
    30.417632891, 30.4176277450001, 30.419248001, 30.4192531460001, 
    30.41979323, 30.4203333140001, 30.4203384590001, 30.4206085000001, 
    30.4206136440001, 30.4203436020001, 30.4203487450001, 30.4200787030001, 
    30.4200838450001, 30.4198138030001, 30.4198240850001, 30.4195540430001, 
    30.4195643200001, 30.4192942780001, 30.417944065, 30.417938926, 
    30.41739884, 30.417393701, 30.4163135260001, 30.416308386, 30.416038342, 
    30.4160332010001, 30.4157631570001, 30.4157580150001, 30.4154879710001, 
    30.4154828280001, 30.4152127840001, 30.4152024960001, 30.409662348, 
    30.4096571790001, 30.409927226, 30.4099220570001, 30.410192104, 
    30.410186933, 30.41045698, 30.4104518080001, 30.4107218550001, 
    30.410716682, 30.411256775, 30.4112516020001, 30.412331785, 30.412326611, 
    30.4125966570001, 30.4125759500001, 30.4128459950001, 30.4128356370001, 
    30.413105682, 30.413100501, 30.4133705460001, 30.4133653640001, 
    30.4136354090001, 30.4136302270001, 30.413900271, 30.4138950880001, 
    30.4141651320001, 30.4141599480001, 30.4144299920001, 30.414424807, 
    30.414694851, 30.414689665, 30.4149597090001, 30.4149545220001, 
    30.4160346960001, 30.4160295080001, 30.4165695940001, 30.4168396370001, 
    30.4168448250001, 30.4171148680001, 30.4171200550001, 30.4173900980001, 
    30.4173952840001, 30.4176653260001, 30.417670512, 30.417940554, 
    30.417950922, 30.4182209640001, 30.4182520470001, 30.4185220890001, 
    30.4185324430001, 30.4188024850001, 30.418812836, 30.4190828770001, 
    30.4190932240001, 30.4193632660001, 30.4193839490001, 30.4196539910001, 
    30.4196849890001, 30.4194149470001, 30.4194768470001, 30.419206805, 
    30.4192119580001, 30.419482, 30.419518043, 30.4197880850001, 30.41979323, 
    30.4192531460001, 30.419248001, 30.4176277450001, 30.417632891, 
    30.4152024960001, 30.4151973510001, 30.414927306, 30.4149118650001, 
    30.4143717760001, 30.414366627, 30.413826537, 30.4138110850001, 
    30.41354104, 30.4135307350001, 30.412990644, 30.41298549, 
    30.4127154440001, 30.412699977, 30.4124299310001, 30.4124247730001, 
    30.412154727, 30.4121444090001, 30.411874363, 30.4118485540001, 
    30.4115785070001, 30.411573343, 30.410763203, 30.410758038, 
    30.4102179440001, 30.410207611, 30.4096675160001, 30.409662348, 
    30.366172625, 30.3661675980001, 30.3664376730001, 30.3664276160001, 
    30.3666976910001, 30.3666825990001, 30.3669526740001, 30.366947641, 
    30.367217716, 30.3672126820001, 30.3677528310001, 30.3677477970001, 
    30.3680178710001, 30.3680027620001, 30.3682728360001, 30.368267798, 
    30.368537872, 30.3685277930001, 30.3687978670001, 30.3687827420001, 
    30.3690528160001, 30.369037683, 30.3698479020001, 30.369852947, 
    30.371473381, 30.3714784250001, 30.372828783, 30.3728237380001, 
    30.373633951, 30.3736389950001, 30.3739090660001, 30.373919152, 
    30.374189222, 30.374199305, 30.374469375, 30.3744744150001, 
    30.3747444850001, 30.374749524, 30.375019594, 30.3750246330001, 
    30.3752947020001, 30.3752997400001, 30.3755698100001, 30.3755748460001, 
    30.3758449160001, 30.3758499510001, 30.376660159, 30.3766651940001, 
    30.3774754, 30.3774804340001, 30.378020571, 30.3780256040001, 
    30.3788358080001, 30.3788408400001, 30.379651043, 30.379656074, 
    30.379926142, 30.3799311720001, 30.3804713060001, 30.380481365, 
    30.3807514310001, 30.3807564590001, 30.381026526, 30.3810214980001, 
    30.381291565, 30.3812865360001, 30.381826668, 30.3818216380001, 
    30.38236177, 30.382631836, 30.382626805, 30.3828968710001, 
    30.3829019020001, 30.3839821620001, 30.3839871920001, 30.3847973860001, 
    30.384802415, 30.3861527350001, 30.386157763, 30.3866978900001, 
    30.386702917, 30.3891334800001, 30.389138507, 30.3899486920001, 
    30.389943665, 30.3902137270001, 30.390208699, 30.3904787600001, 
    30.390473732, 30.392364156, 30.392359126, 30.3928992460001, 30.392904275, 
    30.393174335, 30.3931793630001, 30.3934494230001, 30.39345445, 
    30.39372451, 30.3937295370001, 30.3939995960001, 30.3940046220001, 
    30.395354915, 30.39535994, 30.3959000560001, 30.395905081, 30.396175139, 
    30.396185184, 30.3964552420001, 30.396460264, 30.3980806070001, 
    30.3980755860001, 30.3996959240001, 30.3997009450001, 30.4002410570001, 
    30.4002460780001, 30.4013262990001, 30.4013212780001, 30.402131442, 
    30.4021264200001, 30.4026665280001, 30.4026615060001, 30.4034716670001, 
    30.4034666430001, 30.4042768040001, 30.4042717790001, 30.406972302, 
    30.406967277, 30.4077774310001, 30.4077824560001, 30.4083225580001, 
    30.4083275830001, 30.408597634, 30.4086026580001, 30.408872708, 
    30.4088777310001, 30.409147782, 30.409152804, 30.4102330040001, 
    30.410227982, 30.4110381300001, 30.411033107, 30.4118432540001, 
    30.4118382300001, 30.4123783270001, 30.412373302, 30.4134534940001, 
    30.4134484680001, 30.4139885640001, 30.413983537, 30.4145236310001, 
    30.4145186040001, 30.4150586970001, 30.415063725, 30.415873865, 
    30.4158688370001, 30.41640893, 30.416403901, 30.4172140380001, 
    30.417209008, 30.417749099, 30.4177541290001, 30.4193743970001, 
    30.4193693670001, 30.419639412, 30.419634381, 30.419904425, 30.419899393, 
    30.420169437, 30.420164405, 30.420704492, 30.4206994580001, 30.421509588, 
    30.421504553, 30.422584724, 30.422579689, 30.422849731, 30.422844695, 
    30.423114737, 30.4231097000001, 30.4233797410001, 30.423374703, 
    30.423644745, 30.4236397060001, 30.423909748, 30.4239047080001, 
    30.424174749, 30.4241697080001, 30.42443975, 30.4247097910001, 
    30.4247148310001, 30.424984872, 30.4249899120001, 30.4252599530001, 
    30.4252750680001, 30.4255451080001, 30.425550145, 30.4258201850001, 
    30.425825221, 30.4260952610001, 30.4261002960001, 30.426370336, 
    30.4263753700001, 30.42664541, 30.426650443, 30.4269204830001, 
    30.4269255150001, 30.4274655940001, 30.4274706250001, 30.427740665, 
    30.4277456950001, 30.428015734, 30.4280207640001, 30.4288308810001, 
    30.428835909, 30.4293759870001, 30.429381015, 30.429651053, 30.42965608, 
    30.429926118, 30.4299311440001, 30.4302011820001, 30.430206207, 
    30.4307462830001, 30.430751307, 30.431021345, 30.4310263680001, 
    30.4312964060001, 30.431301429, 30.431571466, 30.4315764880001, 
    30.432116562, 30.432121583, 30.432661657, 30.4326716950001, 
    30.4324016590001, 30.4324066770001, 30.4321366400001, 30.432146673, 
    30.431876636, 30.431886666, 30.431616628, 30.431621642, 30.431351604, 
    30.431361629, 30.431091591, 30.4311016120001, 30.430831574, 30.430836583, 
    30.430566545, 30.4305765600001, 30.430306522, 30.430316534, 30.430046496, 
    30.430056504, 30.4297864650001, 30.42979647, 30.4295264310001, 
    30.429531432, 30.429261393, 30.4292713930001, 30.429001353, 
    30.4290113490001, 30.4287413100001, 30.4287463060001, 30.4284762670001, 
    30.428486257, 30.4282162170001, 30.4282262040001, 30.4279561640001, 
    30.427961156, 30.4276911160001, 30.4277010980001, 30.427431057, 
    30.4274410350001, 30.427170995, 30.4271759820001, 30.4269059420001, 
    30.4269159140001, 30.426645873, 30.4266558420001, 30.426385801, 
    30.426395767, 30.4261257250001, 30.426130707, 30.4258606650001, 
    30.4258706250001, 30.4256005840001, 30.42561054, 30.425340498, 
    30.425345475, 30.4250754330001, 30.425080409, 30.4248103670001, 
    30.424820316, 30.4245502740001, 30.42456022, 30.424290177, 30.424295149, 
    30.424025106, 30.424035046, 30.42349496, 30.4234999290001, 
    30.4229598430001, 30.422964811, 30.4226947670001, 30.422699734, 
    30.4221596470001, 30.4221646130001, 30.421624525, 30.42162949, 
    30.420009222, 30.4200141860001, 30.418123866, 30.4181288290001, 
    30.4165085490001, 30.4165135110001, 30.415433321, 30.415438282, 
    30.4146281380001, 30.414633098, 30.413552904, 30.413547943, 30.413277894, 
    30.413282855, 30.4116625570001, 30.4116675160001, 30.4111274160001, 
    30.411132374, 30.409242018, 30.4092370600001, 30.408156852, 30.408151893, 
    30.407341736, 30.4073367760001, 30.4070667240001, 30.4070716840001, 
    30.4068016310001, 30.4067966710001, 30.405716458, 30.4057114980001, 
    30.4049013370001, 30.4048963750001, 30.404356267, 30.404351304, 
    30.403811196, 30.4038062320001, 30.403266123, 30.4032611590001, 
    30.402721049, 30.4027160840001, 30.4021759730001, 30.402171007, 
    30.401630896, 30.401625929, 30.401355874, 30.4013509060001, 
    30.4008107940001, 30.4008058250001, 30.4002657130001, 30.400260743, 
    30.3999906870001, 30.3999857170001, 30.39971566, 30.3997106890001, 
    30.3994406320001, 30.3994356600001, 30.3972752, 30.397280172, 
    30.3967400550001, 30.3967450260001, 30.3962049080001, 30.396209879, 
    30.39593982, 30.3959447890001, 30.3954046700001, 30.395409639, 
    30.395139579, 30.395144546, 30.394874487, 30.394879453, 30.394609394, 
    30.3946143590001, 30.3940742390001, 30.394079204, 30.3938091430001, 
    30.393814107, 30.393544047, 30.393549009, 30.393278949, 30.393283911, 
    30.3927437890001, 30.3927487500001, 30.392478689, 30.392483649, 
    30.391943526, 30.3919385660001, 30.391668505, 30.391663544, 30.39112342, 
    30.3911184580001, 30.3900382090001, 30.3900431710001, 30.3895030460001, 
    30.389508006, 30.388697817, 30.388692856, 30.3881527290001, 
    30.3881477680001, 30.3878777040001, 30.387872741, 30.3873326140001, 
    30.38732765, 30.386517457, 30.3865124930001, 30.3851621680001, 
    30.3851572030001, 30.384347006, 30.384342041, 30.384071975, 30.384067008, 
    30.3837969420001, 30.3837919740001, 30.383521908, 30.3835169400001, 
    30.3832468730001, 30.383241904, 30.3829718370001, 30.3829668670001, 
    30.382426734, 30.382421763, 30.3821516960001, 30.3821467240001, 
    30.3818766570001, 30.381871684, 30.381331549, 30.381326576, 30.381056508, 
    30.3810515340001, 30.380781466, 30.3807764900001, 30.380506423, 
    30.380501446, 30.3802313780001, 30.3802264010001, 30.3799563330001, 
    30.3799513550001, 30.379681287, 30.3796663470001, 30.379396279, 
    30.379381331, 30.379111263, 30.3790963070001, 30.378826239, 30.378821252, 
    30.3785511830001, 30.3785461950001, 30.378006058, 30.378001069, 
    30.377731, 30.3777260100001, 30.3771858710001, 30.3771808810001, 
    30.3769108120001, 30.37690582, 30.376365681, 30.376360688, 30.376090618, 
    30.376085625, 30.375545485, 30.375540491, 30.375270421, 30.3752654260001, 
    30.3749953550001, 30.37499036, 30.374720289, 30.374705297, 
    30.3744352260001, 30.374425226, 30.374155155, 30.3741501550001, 
    30.3738800830001, 30.373870079, 30.373600008, 30.373595004, 30.373324933, 
    30.3733199280001, 30.3730498570001, 30.373044851, 30.3719645630001, 
    30.371969569, 30.3708892780001, 30.3708842730001, 30.3703441270001, 
    30.370339121, 30.369798974, 30.3697939670001, 30.3695238940001, 
    30.369513877, 30.3692438030001, 30.3692387940001, 30.3689687200001, 
    30.3689637100001, 30.368693636, 30.368683612, 30.368413538, 
    30.3683934800001, 30.3681234060001, 30.368088271, 30.3678181970001, 
    30.367813174, 30.3675431, 30.3675380760001, 30.3672680010001, 
    30.3672629770001, 30.3669929020001, 30.366987877, 30.366177651, 
    30.366172625, 30.390948403, 30.390943362, 30.3912134230001, 
    30.3911932500001, 30.3914633110001, 30.391458265, 30.3917283260001, 
    30.3917232790001, 30.3930735770001, 30.3930786240001, 30.3938888010001, 
    30.393893846, 30.394433963, 30.3944390080001, 30.3974096420001, 
    30.397404597, 30.39929499, 30.3992899450001, 30.400100111, 30.400095064, 
    30.401445338, 30.40144029, 30.403060613, 30.403065661, 30.4054961360001, 
    30.4054910880001, 30.407381448, 30.407376399, 30.408186551, 
    30.4081815010001, 30.4087216020001, 30.4087165510001, 30.410336849, 
    30.4103418990001, 30.411152046, 30.411146995, 30.4114170440001, 
    30.4114119920001, 30.4116820400001, 30.411671934, 30.4119419830001, 
    30.411936928, 30.4124770240001, 30.412471969, 30.412742017, 
    30.4127369600001, 30.4130070080001, 30.4130019510001, 30.413271998, 
    30.41326694, 30.415697359, 30.415702418, 30.416242509, 30.416247566, 
    30.4165176120001, 30.4165125540001, 30.4167826, 30.416777542, 
    30.4170475870001, 30.417042528, 30.417852662, 30.4178577210001, 
    30.41839781, 30.418402869, 30.4194830450001, 30.4194779860001, 
    30.4200180730001, 30.420023132, 30.420833261, 30.420838319, 
    30.4221885310001, 30.422193588, 30.4230037140001, 30.42300877, 
    30.4235488530001, 30.4235589620001, 30.423829003, 30.423834056, 
    30.4241040970001, 30.424134398, 30.4244044390001, 30.42443975, 
    30.4241697080001, 30.424174749, 30.4239047080001, 30.423909748, 
    30.4236397060001, 30.423644745, 30.423374703, 30.4233797410001, 
    30.4231097000001, 30.423114737, 30.422844695, 30.422849731, 30.422579689, 
    30.422584724, 30.421504553, 30.421509588, 30.4206994580001, 30.420704492, 
    30.420164405, 30.420169437, 30.419899393, 30.419904425, 30.419634381, 
    30.419639412, 30.4193693670001, 30.4193743970001, 30.4177541290001, 
    30.417749099, 30.417209008, 30.4172140380001, 30.416403901, 30.41640893, 
    30.4158688370001, 30.415873865, 30.415063725, 30.4150586970001, 
    30.4145186040001, 30.4145236310001, 30.413983537, 30.4139885640001, 
    30.4134484680001, 30.4134534940001, 30.412373302, 30.4123783270001, 
    30.4118382300001, 30.4118432540001, 30.411033107, 30.4110381300001, 
    30.410227982, 30.4102330040001, 30.409152804, 30.409147782, 
    30.4088777310001, 30.408872708, 30.4086026580001, 30.408597634, 
    30.4083275830001, 30.4083225580001, 30.4077824560001, 30.4077774310001, 
    30.406967277, 30.406972302, 30.4042717790001, 30.4042768040001, 
    30.4034666430001, 30.4034716670001, 30.4026615060001, 30.4026665280001, 
    30.4021264200001, 30.402131442, 30.4013212780001, 30.4013262990001, 
    30.4002460780001, 30.4002410570001, 30.3997009450001, 30.3996959240001, 
    30.3980755860001, 30.3980806070001, 30.396460264, 30.3964552420001, 
    30.396185184, 30.396175139, 30.395905081, 30.3959000560001, 30.39535994, 
    30.395354915, 30.3940046220001, 30.3939995960001, 30.3937295370001, 
    30.39372451, 30.39345445, 30.3934494230001, 30.3931793630001, 
    30.393174335, 30.392904275, 30.3928992460001, 30.3928891840001, 
    30.3926191250001, 30.3926040260001, 30.392333966, 30.3923289310001, 
    30.3920588710001, 30.3920538360001, 30.3917837760001, 30.391773702, 
    30.391503642, 30.3914986030001, 30.3912285430001, 30.3912184640001, 
    30.390948403, 30.4192942780001, 30.4195643200001, 30.4195540430001, 
    30.4198240850001, 30.4198138030001, 30.4200838450001, 30.4200787030001, 
    30.4203487450001, 30.4203436020001, 30.4206136440001, 30.4206085000001, 
    30.42059821, 30.421138292, 30.4211279990001, 30.4208579570001, 
    30.42084766, 30.4211177010001, 30.4211074, 30.4213774410001, 
    30.4213619830001, 30.4216320240001, 30.421621714, 30.421891755, 
    30.4218865980001, 30.422156639, 30.4221514820001, 30.422421522, 
    30.4224163640001, 30.422686404, 30.422681245, 30.4229512850001, 
    30.4229306400001, 30.42320068, 30.4231903520001, 30.423460391, 
    30.4234345560001, 30.4237045950001, 30.423678738, 30.423408699, 
    30.423372461, 30.4236425010001, 30.423580278, 30.423310239, 
    30.4232790790001, 30.423549118, 30.423533526, 30.423263488, 
    30.4232530890001, 30.42298305, 30.422972648, 30.4227026090001, 
    30.422681793, 30.422951832, 30.422936211, 30.4232062500001, 30.423201041, 
    30.4234710800001, 30.423455448, 30.423725486, 30.4237098470001, 
    30.4239798850001, 30.4239642370001, 30.4242342750001, 30.424208177, 
    30.4244782150001, 30.424462546, 30.424732583, 30.424727359, 30.424997396, 
    30.424976488, 30.425246525, 30.4252099010001, 30.425479938, 30.425474702, 
    30.4260147750001, 30.4260095390001, 30.426279575, 30.426274338, 
    30.4265443740001, 30.426539136, 30.4270792080001, 30.427084446, 
    30.427894553, 30.4278997910001, 30.428709896, 30.428715133, 
    30.4295252370001, 30.4295304730001, 30.430610609, 30.430615844, 
    30.4314259450001, 30.4314311790001, 30.432241279, 30.4322465120001, 
    30.4330566100001, 30.4330618430001, 30.4333318750001, 30.4333371070001, 
    30.4336071390001, 30.433601907, 30.4338719400001, 30.4338771710001, 
    30.4341472030001, 30.4341524340001, 30.4344224660001, 30.4344276950001, 
    30.4346977270001, 30.434702956, 30.434972988, 30.434978216, 
    30.4355182780001, 30.435523506, 30.4363335990001, 30.4363388250001, 
    30.436878886, 30.436884112, 30.4371541420001, 30.437159367, 
    30.4374293970001, 30.43743462, 30.437704651, 30.4377098730001, 
    30.437979903, 30.4379851250001, 30.438255155, 30.4382708160001, 
    30.438540846, 30.438551282, 30.438821311, 30.4388369590001, 30.439106988, 
    30.4391226280001, 30.439392657, 30.4393978680001, 30.439667898, 
    30.4396783180001, 30.439948347, 30.439953556, 30.440223584, 30.440228792, 
    30.4404988210001, 30.4405040280001, 30.4407740570001, 30.440779263, 
    30.4421294040001, 30.4421346090001, 30.443484746, 30.4434899510001, 
    30.44511011, 30.4451153140001, 30.451595895, 30.451601098, 
    30.4518711200001, 30.4518763230001, 30.4521463450001, 30.452151546, 
    30.452421568, 30.452431968, 30.45270199, 30.452707189, 30.4529772110001, 
    30.4529824090001, 30.4532524300001, 30.453257627, 30.4535276490001, 
    30.453532845, 30.453802866, 30.4538080610001, 30.454078082, 
    30.4540832770001, 30.4543532980001, 30.4543584910001, 30.4546285120001, 
    30.454633705, 30.4549037260001, 30.454914108, 30.455184129, 30.455194508, 
    30.4554645280001, 30.455469717, 30.455739737, 30.455744924, 30.456014945, 
    30.4560201310001, 30.4560253170001, 30.455485276, 30.4554904610001, 
    30.4552204400001, 30.455225624, 30.454955603, 30.4549607860001, 
    30.4546907650001, 30.4546959470001, 30.4544259260001, 30.4544311070001, 
    30.4541610860001, 30.4541662660001, 30.4538962450001, 30.4539066020001, 
    30.4536365810001, 30.4536417580001, 30.4533717370001, 30.4533872640001, 
    30.4531172420001, 30.453127588, 30.452857566, 30.4528627380001, 
    30.452592716, 30.452608227, 30.4523382040001, 30.452353707, 30.452083685, 
    30.4520991790001, 30.4518291570001, 30.45183432, 30.4515642970001, 
    30.451569459, 30.451029412, 30.4510345730001, 30.4504945260001, 
    30.450499687, 30.4502296630001, 30.450234822, 30.4496947740001, 
    30.449699932, 30.4494299080001, 30.449435066, 30.4488950160001, 
    30.448900173, 30.4486301480001, 30.448635304, 30.448365279, 30.448370434, 
    30.447830384, 30.447835538, 30.447565512, 30.4475706650001, 30.447300639, 
    30.4473057920001, 30.4470357660001, 30.447040917, 30.446770891, 
    30.4467811910001, 30.4465111650001, 30.4465163130001, 30.4462462870001, 
    30.4462514350001, 30.4459814080001, 30.445986555, 30.445716528, 
    30.445721674, 30.445451647, 30.4454567920001, 30.4449167380001, 
    30.444927025, 30.444656998, 30.44466214, 30.4443921120001, 30.444397254, 
    30.444127226, 30.4441323660001, 30.4438623390001, 30.4438674780001, 
    30.44359745, 30.4436025890001, 30.44333256, 30.4433376980001, 
    30.442797641, 30.442802778, 30.4419926910001, 30.4419978270001, 
    30.440377649, 30.4403827840001, 30.439842723, 30.4398478580001, 
    30.4374175770001, 30.4374227100001, 30.4366126140001, 30.436617746, 
    30.436077681, 30.4360828120001, 30.4352727130001, 30.4352778430001, 
    30.434467743, 30.4344626130001, 30.4333824770001, 30.433377346, 
    30.432837277, 30.4328321450001, 30.4309418990001, 30.4309470310001, 
    30.429326814, 30.4293319450001, 30.428521835, 30.4285269650001, 
    30.427716853, 30.4277117230001, 30.426361533, 30.4263564020001, 
    30.4250062090001, 30.425011339, 30.4236611420001, 30.4236662710001, 
    30.4228561510001, 30.4228612800001, 30.422051158, 30.4220460290001, 
    30.4215059470001, 30.421500817, 30.4212307760001, 30.421225646, 
    30.420955604, 30.4209504730001, 30.4206804310001, 30.420675299, 
    30.4204052580001, 30.4204001250001, 30.4201300830001, 30.4201249490001, 
    30.4198549070001, 30.4198446360001, 30.419574594, 30.4195694580001, 
    30.4192994150001, 30.4192942780001, 30.410449193, 30.4107192380001, 
    30.4107245020001, 30.410994546, 30.4109998100001, 30.411809943, 
    30.411815205, 30.4128953810001, 30.4128901190001, 30.413430206, 
    30.4134249420001, 30.4139650280001, 30.413959764, 30.41449985, 
    30.414769892, 30.4147751570001, 30.4150451990001, 30.4150557250001, 
    30.4153257670001, 30.4153310290001, 30.415601071, 30.415606332, 
    30.4158763740001, 30.4158816340001, 30.416151676, 30.416162193, 
    30.4164322350001, 30.4164374920001, 30.4167075340001, 30.416718046, 
    30.4169880870001, 30.417014352, 30.417284393, 30.4172948930001, 
    30.417564934, 30.4175754300001, 30.4178454710001, 30.4178507180001, 
    30.4183908000001, 30.4183960460001, 30.418666086, 30.418671331, 
    30.4189413720001, 30.418946616, 30.4192166560001, 30.4192219, 
    30.41976198, 30.4197672220001, 30.4205773420001, 30.4205825830001, 
    30.4211226620001, 30.4211279030001, 30.422208058, 30.422213298, 
    30.4230234140001, 30.4230286530001, 30.4235687290001, 30.423573967, 
    30.423844005, 30.4238492420001, 30.4241192800001, 30.4241245160001, 
    30.4246645910001, 30.4246698260001, 30.4252099010001, 30.425246525, 
    30.424976488, 30.424997396, 30.424727359, 30.424732583, 30.424462546, 
    30.4244782150001, 30.424208177, 30.4242342750001, 30.4239642370001, 
    30.4239798850001, 30.4237098470001, 30.423725486, 30.423455448, 
    30.4234710800001, 30.423201041, 30.4232062500001, 30.422936211, 
    30.422951832, 30.422681793, 30.4227026090001, 30.422972648, 30.42298305, 
    30.4232530890001, 30.423263488, 30.423533526, 30.423549118, 
    30.4232790790001, 30.423310239, 30.423580278, 30.4236425010001, 
    30.423372461, 30.423408699, 30.423678738, 30.4237045950001, 
    30.4234345560001, 30.423460391, 30.4231903520001, 30.42320068, 
    30.4229306400001, 30.4229512850001, 30.422681245, 30.422686404, 
    30.4224163640001, 30.422421522, 30.4221514820001, 30.422156639, 
    30.4218865980001, 30.421891755, 30.421621714, 30.4216320240001, 
    30.4213619830001, 30.4213774410001, 30.4211074, 30.4211177010001, 
    30.42084766, 30.4208579570001, 30.4211279990001, 30.421138292, 
    30.42059821, 30.4206085000001, 30.4203384590001, 30.4203333140001, 
    30.41979323, 30.4197880850001, 30.419518043, 30.419482, 30.4192119580001, 
    30.419206805, 30.4194768470001, 30.4194149470001, 30.4196849890001, 
    30.4196539910001, 30.4193839490001, 30.4193632660001, 30.4190932240001, 
    30.4190828770001, 30.418812836, 30.4188024850001, 30.4185324430001, 
    30.4185220890001, 30.4182520470001, 30.4182209640001, 30.417950922, 
    30.417940554, 30.417670512, 30.4176653260001, 30.4173952840001, 
    30.4173900980001, 30.4171200550001, 30.4171148680001, 30.4168448250001, 
    30.4168396370001, 30.4165695940001, 30.4165124680001, 30.4162424250001, 
    30.416169563, 30.415899521, 30.4158943090001, 30.4156242670001, 
    30.415619055, 30.415349012, 30.415338585, 30.415068542, 30.415063327, 
    30.414793284, 30.4147880680001, 30.4145180250001, 30.414512809, 
    30.414242765, 30.4142375480001, 30.4142323300001, 30.4139622860001, 
    30.4139518470001, 30.413681803, 30.4136713610001, 30.413401317, 
    30.4133960940001, 30.4131260500001, 30.4131208270001, 30.4128507830001, 
    30.4128455580001, 30.412575514, 30.412570289, 30.4123002440001, 
    30.4122950180001, 30.412024973, 30.412014519, 30.411744474, 30.411734016, 
    30.411463971, 30.4114587400001, 30.4111886950001, 30.4111677650001, 
    30.41089772, 30.4108767750001, 30.41060673, 30.4105805290001, 
    30.410310484, 30.4102842610001, 30.410014215, 30.4100089680001, 
    30.410279014, 30.410221236, 30.4099511900001, 30.4099354140001, 
    30.4102054590001, 30.410200199, 30.4104702440001, 30.410449193, 
    30.3943565530001, 30.394330317, 30.394600371, 30.3945951210001, 
    30.3948651760001, 30.394859925, 30.395129979, 30.3951247270001, 
    30.395664835, 30.395654329, 30.3959243830001, 30.3959191280001, 
    30.3961891820001, 30.39617867, 30.396448724, 30.3964434660001, 
    30.3969835730001, 30.396978314, 30.397248367, 30.3972431080001, 
    30.3975131610001, 30.397507901, 30.397777954, 30.397772693, 
    30.3980427450001, 30.3980374830001, 30.3983075360001, 30.3983022730001, 
    30.398572325, 30.398551266, 30.3988213170001, 30.3988160500001, 
    30.3985459990001, 30.398540731, 30.3988107820001, 30.3988055140001, 
    30.399075565, 30.3990702950001, 30.3993403470001, 30.3993350760001, 
    30.399605127, 30.3996103980001, 30.4006906010001, 30.400695871, 
    30.4012359720001, 30.401241241, 30.402321441, 30.4023267090001, 
    30.4028668080001, 30.4028720750001, 30.403952271, 30.403947004, 
    30.406647483, 30.406642215, 30.4085325400001, 30.4085378090001, 
    30.4088078550001, 30.408813122, 30.4093532140001, 30.409358481, 
    30.409898571, 30.4099038370001, 30.4104439280001, 30.410449193, 
    30.4104702440001, 30.410200199, 30.4102054590001, 30.4099354140001, 
    30.4099511900001, 30.410221236, 30.410279014, 30.4100089680001, 
    30.410014215, 30.4102842610001, 30.410310484, 30.4105805290001, 
    30.41060673, 30.4108767750001, 30.41089772, 30.4111677650001, 
    30.4111886950001, 30.4114587400001, 30.411463971, 30.411734016, 
    30.411744474, 30.412014519, 30.412024973, 30.4122950180001, 
    30.4123002440001, 30.412570289, 30.412575514, 30.4128455580001, 
    30.4128507830001, 30.4131208270001, 30.4131260500001, 30.4133960940001, 
    30.413401317, 30.4136713610001, 30.413681803, 30.4139518470001, 
    30.4139622860001, 30.4142323300001, 30.4142375480001, 30.4128873270001, 
    30.412892544, 30.4126225000001, 30.412627716, 30.4123576710001, 
    30.412368101, 30.412098056, 30.41210327, 30.4112931340001, 
    30.4112879210001, 30.411017875, 30.411023088, 30.4102129510001, 
    30.410218163, 30.407247646, 30.4067075500001, 30.4067023380001, 
    30.4061622410001, 30.4061570280001, 30.40588698, 30.4058817660001, 
    30.4056117170001, 30.405601286, 30.405331237, 30.4053260200001, 
    30.404785922, 30.4047754860001, 30.4045054370001, 30.4045002180001, 
    30.404230168, 30.404224948, 30.4036848490001, 30.4036796280001, 
    30.403409578, 30.4034043560001, 30.402864256, 30.402859033, 
    30.4023189320001, 30.4023137090001, 30.402043658, 30.4020384340001, 
    30.401768383, 30.4017631570001, 30.4014931070001, 30.40148788, 
    30.400947778, 30.4009425510001, 30.4006725, 30.4006672720001, 
    30.4003972200001, 30.400391991, 30.3998518880001, 30.3998466580001, 
    30.399576606, 30.399560912, 30.3992908600001, 30.3992856260001, 
    30.399015574, 30.3990103400001, 30.398470235, 30.398465, 
    30.3979248950001, 30.397903946, 30.397633893, 30.3976286540001, 
    30.3973586010001, 30.3973481190001, 30.3970780660001, 30.3970728240001, 
    30.3968027710001, 30.396797528, 30.395987367, 30.3959821230001, 
    30.3957120690001, 30.395706825, 30.3943565530001, 30.3712653170001, 
    30.372075528, 30.3720703990001, 30.3723404690001, 30.3723353390001, 
    30.3726054090001, 30.3726002780001, 30.3728703470001, 30.372865216, 
    30.373135285, 30.373130153, 30.3736702910001, 30.3736651580001, 
    30.374475364, 30.3744702290001, 30.3747402980001, 30.3747094730001, 
    30.3749795410001, 30.374964117, 30.3752341850001, 30.3752084600001, 
    30.375478528, 30.3754682320001, 30.375738299, 30.37573315, 
    30.3760032170001, 30.375992916, 30.3762629830001, 30.3762423690001, 
    30.375972302, 30.3759619900001, 30.376232057, 30.3762268990001, 
    30.376496966, 30.3764866490001, 30.376216582, 30.3762062610001, 
    30.3759361940001, 30.375931032, 30.3756609650001, 30.3756454740001, 
    30.375915541, 30.375910375, 30.3761804420001, 30.376170109, 
    30.3764401760001, 30.3764350070001, 30.376705074, 30.3766947350001, 
    30.376964801, 30.376959631, 30.3772296970001, 30.377224525, 
    30.3774945910001, 30.377489418, 30.3780295500001, 30.3780192020001, 
    30.377749136, 30.3777439610001, 30.377473895, 30.377463542, 
    30.3771934760001, 30.3771312820001, 30.377401348, 30.3773961590001, 
    30.377666225, 30.3776610350001, 30.3779311010001, 30.37792591, 
    30.378466041, 30.3784608490001, 30.3787309140001, 30.3787257220001, 
    30.3795359160001, 30.379530722, 30.380340915, 30.3803357210001, 
    30.3806057840001, 30.380600589, 30.380870653, 30.380865457, 30.38113552, 
    30.381130324, 30.381400387, 30.381395189, 30.3816652520001, 30.381654854, 
    30.3821949800001, 30.382189779, 30.3824598420001, 30.382449438, 
    30.3827195010001, 30.3827142980001, 30.38298436, 30.3829739510001, 
    30.383244013, 30.3832336, 30.3835036620001, 30.3834932460001, 
    30.383763308, 30.3837528880001, 30.38402295, 30.384012526, 
    30.3845526490001, 30.384547436, 30.384817497, 30.384812283, 
    30.3853524040001, 30.3853471890001, 30.3856172500001, 30.3856120340001, 
    30.386422214, 30.3864169980001, 30.3869571170001, 30.3869519, 
    30.387221959, 30.387216741, 30.387756859, 30.38775164, 30.388021699, 
    30.3880164780001, 30.3882865370001, 30.3882813160001, 30.3885513750001, 
    30.3885461520001, 30.389356327, 30.3893511040001, 30.389621162, 
    30.3896159380001, 30.3904261110001, 30.3904313350001, 30.390701393, 
    30.3907170590001, 30.3909871160001, 30.3910027750001, 30.391272832, 
    30.391288483, 30.3915585400001, 30.3915637550001, 30.3918338120001, 
    30.391849452, 30.3921195080001, 30.39214035, 30.3924104060001, 
    30.3924156140001, 30.392685671, 30.3926908780001, 30.392960934, 
    30.392966141, 30.3932361970001, 30.3932414020001, 30.393511458, 
    30.3935166630001, 30.394056774, 30.394061978, 30.394602089, 30.394607292, 
    30.394877347, 30.394882549, 30.395152604, 30.395157806, 30.395697915, 
    30.3957031160001, 30.396243225, 30.3962484240001, 30.3967885330001, 
    30.3967937310001, 30.397063786, 30.3970741800001, 30.3973442340001, 
    30.397354625, 30.397624679, 30.397629873, 30.397899927, 30.3979051200001, 
    30.398175173, 30.398185557, 30.398455611, 30.398465991, 30.398736044, 
    30.3987412330001, 30.399551392, 30.39955658, 30.4003667380001, 
    30.4003719250001, 30.400912029, 30.400917216, 30.4011872670001, 
    30.4011924530001, 30.401462505, 30.4014676890001, 30.401737741, 
    30.4017429250001, 30.402012976, 30.4020181590001, 30.4022882100001, 
    30.4022985730001, 30.402568624, 30.4025945160001, 30.4028645670001, 
    30.4028852650001, 30.403155316, 30.4031656600001, 30.4034357100001, 
    30.403461554, 30.403731604, 30.40373677, 30.4040068210001, 
    30.4040119860001, 30.404282037, 30.404287201, 30.404557251, 30.4045779, 
    30.4043078490001, 30.4043336390001, 30.404063588, 30.404073898, 
    30.403533796, 30.40353895, 30.4032688990001, 30.4032843540001, 
    30.403014302, 30.403019452, 30.4027494010001, 30.4027545500001, 
    30.402484498, 30.402489646, 30.402219594, 30.4022247410001, 30.401954689, 
    30.4019598360001, 30.4016897830001, 30.401694929, 30.4011548240001, 
    30.4011599680001, 30.4008899150001, 30.4008950590001, 30.400625006, 
    30.4006301490001, 30.400360096, 30.400370378, 30.400100325, 30.400105465, 
    30.3998354120001, 30.3998405510001, 30.3995704970001, 30.3995756350001, 
    30.3993055820001, 30.399310719, 30.399040665, 30.399050937, 30.398780883, 
    30.3987860170001, 30.3985159630001, 30.398526229, 30.398256175, 
    30.398261307, 30.3979912520001, 30.3979963830001, 30.397726328, 
    30.3977314580001, 30.3974614030001, 30.3974767880001, 30.3972067330001, 
    30.39722211, 30.396952055, 30.396962301, 30.396692246, 30.3967024890001, 
    30.3961623770001, 30.3961674970001, 30.3956273850001, 30.395632504, 
    30.395092391, 30.39509751, 30.3948274530001, 30.394557396, 30.394552278, 
    30.394282221, 30.3942771010001, 30.394007044, 30.3940019240001, 
    30.3937318660001, 30.393726745, 30.3934566880001, 30.3934515660001, 
    30.3931815080001, 30.3931763860001, 30.392906328, 30.3929012040001, 
    30.3918209710001, 30.391815847, 30.3912757300001, 30.3912808540001, 
    30.3904706770001, 30.3904758, 30.390205741, 30.390210864, 30.389940804, 
    30.3899459260001, 30.3896758660001, 30.3896809870001, 30.389410927, 
    30.3894160470001, 30.3888759270001, 30.3888810460001, 30.3886109850001, 
    30.3886212210001, 30.3883511600001, 30.388356276, 30.388086216, 
    30.3880913310001, 30.3878212700001, 30.387831498, 30.3872913760001, 
    30.3873016000001, 30.3870315390001, 30.38703665, 30.3867665880001, 
    30.3867614770001, 30.386491415, 30.3864863040001, 30.386216242, 
    30.3862111290001, 30.3856710050001, 30.385665891, 30.3837754520001, 
    30.3837805650001, 30.382970374, 30.3829754870001, 30.3810850360001, 
    30.3810901470001, 30.380009886, 30.380004775, 30.3773041110001, 
    30.3772989980001, 30.3762187290001, 30.3762238410001, 30.3754136370001, 
    30.3754085240001, 30.3751384560001, 30.3751333430001, 30.3735129300001, 
    30.373507816, 30.3732377470001, 30.3732326320001, 30.3729625620001, 
    30.3729523310001, 30.3726822610001, 30.3726771440001, 30.372407074, 
    30.372401956, 30.372131886, 30.3721062820001, 30.3718362120001, 
    30.3718310880001, 30.3715610180001, 30.3715507680001, 30.3712806980001, 
    30.3712653170001, 30.364360102, 30.3643549010001, 30.364624974, 
    30.364619772, 30.3648898440001, 30.3648846410001, 30.365154714, 
    30.3651443050001, 30.365414377, 30.365403965, 30.3656740370001, 
    30.3656688300001, 30.365938902, 30.3659284840001, 30.3664686270001, 
    30.366463417, 30.3667334890001, 30.3667230660001, 30.3669931370001, 
    30.36697228, 30.3672423510001, 30.3672371340001, 30.367507205, 
    30.3675019880001, 30.3680421290001, 30.368036911, 30.368577052, 
    30.368571832, 30.369111972, 30.3691067520001, 30.3699169610001, 
    30.369922181, 30.3704623200001, 30.3704675390001, 30.3726280870001, 
    30.3726228680001, 30.3731630030001, 30.3731316670001, 30.3734017350001, 
    30.3733912820001, 30.3736613500001, 30.373650894, 30.3739209610001, 
    30.3739157310001, 30.374185798, 30.374154403, 30.3738843370001, 
    30.3738738650001, 30.373603798, 30.3735985610001, 30.3733284940001, 
    30.373318016, 30.3730479490001, 30.3730427090001, 30.372772642, 
    30.37276216, 30.3724920920001, 30.37248685, 30.3722167820001, 
    30.372211539, 30.3724816060001, 30.372471117, 30.3727411840001, 
    30.3727359380001, 30.373546139, 30.3735408920001, 30.3743510910001, 
    30.3743458430001, 30.374885976, 30.3748807270001, 30.375150793, 
    30.3751245350001, 30.3753946000001, 30.3753893460001, 30.3756594110001, 
    30.375643643, 30.375913708, 30.375897932, 30.376167997, 30.3761574750001, 
    30.3764275400001, 30.3764222780001, 30.3766923430001, 30.3766870790001, 
    30.3772272080001, 30.377221944, 30.377492008, 30.3774867430001, 
    30.3796472510001, 30.3796525160001, 30.379922579, 30.3799278430001, 
    30.380197906, 30.380203169, 30.380473232, 30.380478495, 30.3807485570001, 
    30.3807538190001, 30.3812939430001, 30.3812992040001, 30.3834596950001, 
    30.3834649550001, 30.3840050760001, 30.384010335, 30.3842803950001, 
    30.3842856540001, 30.3856359530001, 30.3856412110001, 30.3867214480001, 
    30.3867267040001, 30.3872668220001, 30.3872825870001, 30.387552645, 
    30.3875578980001, 30.3878279570001, 30.3878384600001, 30.3881085190001, 
    30.388119019, 30.3883890770001, 30.388394326, 30.3889344420001, 
    30.388939689, 30.392990539, 30.3929852910001, 30.3937954560001, 
    30.3937902070001, 30.394330317, 30.3943565530001, 30.394086498, 
    30.394091743, 30.3935516330001, 30.393556877, 30.3930167660001, 
    30.393022009, 30.392481897, 30.392487139, 30.392217083, 30.3922275640001, 
    30.3919575080001, 30.391962747, 30.391422634, 30.39143311, 
    30.3911630530001, 30.3911682900001, 30.390898233, 30.3909034690001, 
    30.3906334120001, 30.3906386460001, 30.390368589, 30.390379056, 
    30.3901089980001, 30.390124691, 30.3898546340001, 30.389875546, 
    30.3901456030001, 30.390150829, 30.3904208860001, 30.3904261110001, 
    30.3896159380001, 30.389621162, 30.3893511040001, 30.389356327, 
    30.3885461520001, 30.3885513750001, 30.3882813160001, 30.3882865370001, 
    30.3880164780001, 30.388021699, 30.38775164, 30.387756859, 30.387216741, 
    30.387221959, 30.3869519, 30.3869571170001, 30.3864169980001, 
    30.386422214, 30.3856120340001, 30.3856172500001, 30.3853471890001, 
    30.3853524040001, 30.384812283, 30.384817497, 30.384547436, 
    30.3845526490001, 30.384012526, 30.38402295, 30.3837528880001, 
    30.383763308, 30.3834932460001, 30.3835036620001, 30.3832336, 
    30.383244013, 30.3829739510001, 30.38298436, 30.3827142980001, 
    30.3827195010001, 30.382449438, 30.3824598420001, 30.382189779, 
    30.3821949800001, 30.381654854, 30.3816652520001, 30.381395189, 
    30.381400387, 30.381130324, 30.38113552, 30.380865457, 30.380870653, 
    30.380600589, 30.3806057840001, 30.3803357210001, 30.380340915, 
    30.379530722, 30.3795359160001, 30.3787257220001, 30.3787309140001, 
    30.3784608490001, 30.378466041, 30.37792591, 30.3779311010001, 
    30.3776610350001, 30.377666225, 30.3773961590001, 30.377401348, 
    30.3771312820001, 30.3771934760001, 30.377463542, 30.377473895, 
    30.3777439610001, 30.377749136, 30.3780192020001, 30.3780295500001, 
    30.377489418, 30.3774945910001, 30.377224525, 30.3772296970001, 
    30.376959631, 30.376964801, 30.3766947350001, 30.376705074, 
    30.3764350070001, 30.3764401760001, 30.376170109, 30.3761804420001, 
    30.375910375, 30.375915541, 30.3756454740001, 30.3756609650001, 
    30.375931032, 30.3759361940001, 30.3762062610001, 30.376216582, 
    30.3764866490001, 30.376496966, 30.3762268990001, 30.376232057, 
    30.3759619900001, 30.375972302, 30.3762423690001, 30.3762629830001, 
    30.375992916, 30.3760032170001, 30.37573315, 30.375738299, 
    30.3754682320001, 30.375478528, 30.3752084600001, 30.3752341850001, 
    30.374964117, 30.3749795410001, 30.3747094730001, 30.3747402980001, 
    30.3744702290001, 30.374475364, 30.3736651580001, 30.3736702910001, 
    30.373130153, 30.373135285, 30.372865216, 30.3728703470001, 
    30.3726002780001, 30.3726054090001, 30.3723353390001, 30.3723404690001, 
    30.3720703990001, 30.372075528, 30.3712653170001, 30.3712601880001, 
    30.3709901180001, 30.370984988, 30.370714918, 30.370704656, 
    30.3704345850001, 30.370429453, 30.3701593820001, 30.3701285700001, 
    30.369858499, 30.3698327980001, 30.3695627270001, 30.3695575840001, 
    30.3692875130001, 30.369277224, 30.369007153, 30.368996861, 30.36872679, 
    30.368721642, 30.3681814990001, 30.368176351, 30.367636207, 30.367631058, 
    30.366820841, 30.3668156910001, 30.366005473, 30.366000322, 30.365730249, 
    30.3657096370001, 30.365439564, 30.3654292530001, 30.36515918, 
    30.3651540230001, 30.364883949, 30.3648736330001, 30.3643334860001, 
    30.3643283260001, 30.3637881780001, 30.363783018, 30.363512944, 
    30.3635077820001, 30.363237708, 30.3631912170001, 30.3629211430001, 
    30.362910802, 30.3631808760001, 30.3631757040001, 30.363445778, 
    30.3634354320001, 30.36397558, 30.363970405, 30.3645105520001, 
    30.3644794860001, 30.364209413, 30.364193867, 30.3639237940001, 
    30.363897868, 30.363627794, 30.3636070370001, 30.3638771110001, 
    30.3638719190001, 30.3644120660001, 30.3644068740001, 30.36494702, 
    30.364936632, 30.3646665590001, 30.364635375, 30.3643653030001, 
    30.364360102, 30.405331237, 30.405601286, 30.4056117170001, 
    30.4058817660001, 30.40588698, 30.4061570280001, 30.4061622410001, 
    30.4067023380001, 30.4067075500001, 30.407247646, 30.407252858, 
    30.4077929530001, 30.407798164, 30.4080682110001, 30.408073421, 
    30.40915361, 30.409158819, 30.4096989120001, 30.4097041200001, 
    30.409974166, 30.409979374, 30.410519466, 30.410514259, 30.4124045770001, 
    30.412414991, 30.412685036, 30.4126902420001, 30.41377042, 
    30.4137652140001, 30.4140352580001, 30.414030052, 30.414300096, 
    30.414294888, 30.4145649320001, 30.4145597240001, 30.4148297670001, 
    30.4148245580001, 30.4150946010001, 30.415089391, 30.415359435, 
    30.4153542230001, 30.4156242670001, 30.4158943090001, 30.415899521, 
    30.416169563, 30.4162424250001, 30.4165124680001, 30.4165695940001, 
    30.4160295080001, 30.4160346960001, 30.4149545220001, 30.4149597090001, 
    30.414689665, 30.414694851, 30.414424807, 30.4144299920001, 
    30.4141599480001, 30.4141651320001, 30.4138950880001, 30.413900271, 
    30.4136302270001, 30.4136354090001, 30.4133653640001, 30.4133705460001, 
    30.413100501, 30.413105682, 30.4128356370001, 30.412565591, 30.412570771, 
    30.41203068, 30.4120203200001, 30.411750274, 30.411745092, 
    30.4114750460001, 30.411464681, 30.4111946350001, 30.4111894500001, 
    30.410919404, 30.4109142190001, 30.410644173, 30.4106182350001, 
    30.4103481880001, 30.410322228, 30.410052181, 30.410041791, 
    30.4097717440001, 30.4097665480001, 30.409496501, 30.409491303, 
    30.4092212570001, 30.409210859, 30.408940812, 30.4089356120001, 
    30.4083955180001, 30.4083903170001, 30.4081202690001, 30.408109865, 
    30.407839817, 30.407834614, 30.4075645660001, 30.407559361, 30.407289314, 
    30.4072841080001, 30.4070140600001, 30.407008854, 30.4067388060001, 
    30.4067335990001, 30.4064635510001, 30.4064583430001, 30.4061882940001, 
    30.4061830850001, 30.4059130370001, 30.4059078270001, 30.405637778, 
    30.405632568, 30.4053625190001, 30.405331237, 30.407247646, 30.410218163, 
    30.4102129510001, 30.411023088, 30.411017875, 30.4112879210001, 
    30.4112931340001, 30.41210327, 30.412098056, 30.412368101, 
    30.4123576710001, 30.412627716, 30.4126225000001, 30.412892544, 
    30.4128873270001, 30.4142375480001, 30.414242765, 30.414512809, 
    30.4145180250001, 30.4147880680001, 30.414793284, 30.415063327, 
    30.415068542, 30.415338585, 30.415349012, 30.415619055, 30.4156242670001, 
    30.4153542230001, 30.415359435, 30.415089391, 30.4150946010001, 
    30.4148245580001, 30.4148297670001, 30.4145597240001, 30.4145649320001, 
    30.414294888, 30.414300096, 30.414030052, 30.4140352580001, 
    30.4137652140001, 30.41377042, 30.4126902420001, 30.412685036, 
    30.412414991, 30.4124045770001, 30.410514259, 30.410519466, 30.409979374, 
    30.409974166, 30.4097041200001, 30.4096989120001, 30.409158819, 
    30.40915361, 30.408073421, 30.4080682110001, 30.407798164, 
    30.4077929530001, 30.407252858, 30.407247646, 30.357313597, 30.357303372, 
    30.3575734510001, 30.3575581060001, 30.3578281850001, 30.3578230680001, 
    30.358093147, 30.358088029, 30.3583581080001, 30.358352989, 
    30.3586230670001, 30.358607707, 30.3583376290001, 30.3583325070001, 
    30.358602585, 30.358597462, 30.3588675400001, 30.358841913, 30.35911199, 
    30.359106862, 30.3593769400001, 30.3593718110001, 30.3596418880001, 
    30.359621363, 30.3598914400001, 30.3598863060001, 30.3601563830001, 
    30.360146113, 30.36041619, 30.3604110540001, 30.36068113, 30.360675993, 
    30.3609460700001, 30.3609409320001, 30.3612110080001, 30.3611750170001, 
    30.361164726, 30.361434801, 30.3614296550001, 30.361969806, 30.361964658, 
    30.362234733, 30.362208981, 30.362479056, 30.3624739030001, 30.362743978, 
    30.3627388240001, 30.363008898, 30.362998588, 30.3632686620001, 
    30.363258348, 30.3635284220001, 30.363523263, 30.3637933380001, 
    30.3637881780001, 30.3643283260001, 30.3643334860001, 30.3648736330001, 
    30.364883949, 30.3651540230001, 30.36515918, 30.3654292530001, 
    30.365439564, 30.3657096370001, 30.365730249, 30.366000322, 30.366005473, 
    30.3668156910001, 30.366820841, 30.367631058, 30.367636207, 30.368176351, 
    30.3681814990001, 30.368721642, 30.36872679, 30.368996861, 30.369007153, 
    30.369277224, 30.3692875130001, 30.3695575840001, 30.3695627270001, 
    30.3698327980001, 30.369858499, 30.3701285700001, 30.3701593820001, 
    30.370429453, 30.3704345850001, 30.370704656, 30.370714918, 30.370984988, 
    30.3709901180001, 30.3712601880001, 30.3712653170001, 30.3712806980001, 
    30.3715507680001, 30.3715610180001, 30.3718310880001, 30.3718362120001, 
    30.3721062820001, 30.372131886, 30.372401956, 30.372407074, 
    30.3726771440001, 30.3726822610001, 30.3729523310001, 30.3729625620001, 
    30.3732326320001, 30.3732377470001, 30.373507816, 30.3735129300001, 
    30.3751333430001, 30.3751384560001, 30.3754085240001, 30.3754136370001, 
    30.3762238410001, 30.37624428, 30.3759742120001, 30.3759793200001, 
    30.3740888400001, 30.3740990520001, 30.3738289830001, 30.373834088, 
    30.3732939490001, 30.373299053, 30.372758913, 30.3727640160001, 
    30.3722238760001, 30.3722289780001, 30.370878625, 30.370883726, 
    30.3703435830001, 30.370348683, 30.3689983240001, 30.369003424, 
    30.3681932060001, 30.368198304, 30.367658159, 30.3676632560001, 
    30.367393183, 30.36739828, 30.3671282060001, 30.3671333020001, 
    30.3649727100001, 30.364977804, 30.364437654, 30.364442748, 30.363902598, 
    30.3639076910001, 30.362557312, 30.3625624040001, 30.3614820980001, 
    30.3614871890001, 30.3612171120001, 30.361227291, 30.3609572140001, 
    30.3609623020001, 30.360692225, 30.3606973120001, 30.360427235, 
    30.3604323210001, 30.360162244, 30.360172414, 30.359632258, 30.359627174, 
    30.3593570960001, 30.3593520100001, 30.359081932, 30.3590768460001, 
    30.3585366890001, 30.358531602, 30.3582615230001, 30.3582309810001, 
    30.3579609020001, 30.35792013, 30.358190209, 30.3581646970001, 
    30.357894619, 30.357874194, 30.3576041150001, 30.3575938970001, 
    30.3573238180001, 30.357313597, 30.347157624, 30.3471525310001, 
    30.3474226160001, 30.3474175220001, 30.3476876070001, 30.3476825120001, 
    30.348222682, 30.348217586, 30.349027839, 30.349022742, 30.34956291, 
    30.3498329930001, 30.3498278960001, 30.3500979790001, 30.350092881, 
    30.3503629640001, 30.350357865, 30.350898031, 30.350892931, 
    30.3511630130001, 30.3511579120001, 30.3514279950001, 30.35141779, 
    30.352228037, 30.3522331390001, 30.352773303, 30.3527682000001, 
    30.3530382820001, 30.353033178, 30.3551938250001, 30.3551887200001, 
    30.3554588000001, 30.3554485870001, 30.355988747, 30.35598364, 
    30.3562537190001, 30.3562486110001, 30.35651869, 30.3565135810001, 
    30.3567836600001, 30.3567785500001, 30.3570486290001, 30.3570435180001, 
    30.357313597, 30.3573238180001, 30.3575938970001, 30.3576041150001, 
    30.357874194, 30.357894619, 30.3581646970001, 30.358190209, 30.35792013, 
    30.3579609020001, 30.3582309810001, 30.3582615230001, 30.358281866, 
    30.3580117880001, 30.3580168710001, 30.35828695, 30.3582920330001, 
    30.35883219, 30.3588423530001, 30.3591124320001, 30.3591225910001, 
    30.359392669, 30.359418052, 30.3596881300001, 30.3596932040001, 
    30.3599632830001, 30.359968356, 30.3602384340001, 30.3602435060001, 
    30.3610537390001, 30.36105881, 30.3615989640001, 30.361869042, 
    30.3618741120001, 30.362144189, 30.362149259, 30.362419335, 30.362424404, 
    30.3626944810001, 30.362699548, 30.3629696250001, 30.362974692, 
    30.3632447680001, 30.363249834, 30.3637899870001, 30.3637950520001, 
    30.3643352030001, 30.364340268, 30.364610343, 30.364615407, 30.364885482, 
    30.364890545, 30.365970845, 30.3659759070001, 30.36678613, 
    30.3667911910001, 30.3670612650001, 30.367066326, 30.366796251, 
    30.3668063690001, 30.3665362950001, 30.366546408, 30.3662763340001, 
    30.3662914980001, 30.3665615730001, 30.3665817790001, 30.3668518540001, 
    30.366856903, 30.3673970520001, 30.3674021, 30.3679422480001, 
    30.3679472960001, 30.368487443, 30.3684924900001, 30.3687625640001, 
    30.3687676100001, 30.369037683, 30.3690528160001, 30.3687827420001, 
    30.3687978670001, 30.3685277930001, 30.368537872, 30.368267798, 
    30.3682728360001, 30.3680027620001, 30.3680178710001, 30.3677477970001, 
    30.3677528310001, 30.3672126820001, 30.367217716, 30.366947641, 
    30.3669526740001, 30.3666825990001, 30.3666976910001, 30.3664276160001, 
    30.3664376730001, 30.3661675980001, 30.366172625, 30.365362399, 
    30.3653573720001, 30.364277067, 30.3642720390001, 30.363731886, 
    30.3637268580001, 30.361836317, 30.3618312880001, 30.360210818, 
    30.3602158480001, 30.359945769, 30.3599507980001, 30.359680719, 
    30.3596857470001, 30.3594156680001, 30.35942572, 30.359155641, 
    30.359160666, 30.3588905870001, 30.358895611, 30.358625531, 
    30.3586305540001, 30.358360475, 30.3583654970001, 30.3580954170001, 
    30.3581004380001, 30.3578303580001, 30.357290198, 30.3572851760001, 
    30.3564749340001, 30.3564699120001, 30.355929749, 30.3559247260001, 
    30.3556546450001, 30.3556496210001, 30.3553795390001, 30.3553745140001, 
    30.3551044330001, 30.35509438, 30.354824299, 30.3548092130001, 
    30.3545391320001, 30.3545290700001, 30.354258988, 30.354253956, 
    30.3539838740001, 30.3539788410001, 30.353438677, 30.3534336430001, 
    30.3528934780001, 30.352888443, 30.3520781940001, 30.3520731580001, 
    30.3518030750001, 30.3517980390001, 30.3515279550001, 30.3515229180001, 
    30.3509827510001, 30.3509777130001, 30.3507076290001, 30.35070259, 
    30.350972674, 30.3509625930001, 30.351232677, 30.3512175500001, 
    30.350947466, 30.3509424220001, 30.351212506, 30.3512074610001, 
    30.351477544, 30.3514674510001, 30.351737535, 30.3517274380001, 
    30.351997522, 30.351987421, 30.3522575040001, 30.3522524530001, 
    30.352522536, 30.352517484, 30.3527875660001, 30.352777459, 
    30.3530475420001, 30.3530222580001, 30.352752176, 30.352747116, 
    30.3524770340001, 30.352471973, 30.3522018910001, 30.35219683, 
    30.3519267470001, 30.351891294, 30.3516212110001, 30.3516110740001, 
    30.351340991, 30.351325778, 30.3510556950001, 30.3510506220001, 
    30.350780539, 30.350770391, 30.3505003080001, 30.350449515, 
    30.3501794320001, 30.3501743480001, 30.349904264, 30.349899179, 
    30.3496290950001, 30.3496240100001, 30.349083842, 30.3490787550001, 
    30.348808671, 30.3488035830001, 30.348533499, 30.34852841, 
    30.3482583260001, 30.3482532360001, 30.347983152, 30.347978062, 
    30.347707977, 30.347702886, 30.3471627160001, 30.347157624 ;

 catchments_node_count = 242, 44, 254, 177, 83, 37, 541, 33, 99, 518, 192, 
    325, 215, 179, 360, 356, 117, 59, 182, 262 ;

 catchments_part_node_count = 242, 44, 254, 177, 5, 78, 37, 541, 33, 99, 518, 
    192, 325, 215, 179, 360, 356, 117, 59, 182, 262 ;

 catchments_AreaSqKM = 3.0861, 0.0738, 4.0752, 2.5803, 0.4923, 0.0801, 
    18.8136, 0.108, 1.0287, 13.3281, 3.006, 9.1854, 3.0861, 2.5344, 8.4861, 
    6.6735, 0.6759, 0.1854, 2.7405, 3.5118 ;
}
